//megafunction wizard: %Altera SOPC Builder%
//GENERATION: STANDARD
//VERSION: WM1.0


//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module button_pio_s1_arbitrator (
                                  // inputs:
                                   button_pio_s1_irq,
                                   button_pio_s1_readdata,
                                   clk,
                                   pb_cpu_to_io_m1_address_to_slave,
                                   pb_cpu_to_io_m1_burstcount,
                                   pb_cpu_to_io_m1_chipselect,
                                   pb_cpu_to_io_m1_latency_counter,
                                   pb_cpu_to_io_m1_read,
                                   pb_cpu_to_io_m1_write,
                                   pb_cpu_to_io_m1_writedata,
                                   reset_n,

                                  // outputs:
                                   button_pio_s1_address,
                                   button_pio_s1_chipselect,
                                   button_pio_s1_irq_from_sa,
                                   button_pio_s1_readdata_from_sa,
                                   button_pio_s1_reset_n,
                                   button_pio_s1_write_n,
                                   button_pio_s1_writedata,
                                   d1_button_pio_s1_end_xfer,
                                   pb_cpu_to_io_m1_granted_button_pio_s1,
                                   pb_cpu_to_io_m1_qualified_request_button_pio_s1,
                                   pb_cpu_to_io_m1_read_data_valid_button_pio_s1,
                                   pb_cpu_to_io_m1_requests_button_pio_s1
                                )
;

  output  [  1: 0] button_pio_s1_address;
  output           button_pio_s1_chipselect;
  output           button_pio_s1_irq_from_sa;
  output  [  2: 0] button_pio_s1_readdata_from_sa;
  output           button_pio_s1_reset_n;
  output           button_pio_s1_write_n;
  output  [  2: 0] button_pio_s1_writedata;
  output           d1_button_pio_s1_end_xfer;
  output           pb_cpu_to_io_m1_granted_button_pio_s1;
  output           pb_cpu_to_io_m1_qualified_request_button_pio_s1;
  output           pb_cpu_to_io_m1_read_data_valid_button_pio_s1;
  output           pb_cpu_to_io_m1_requests_button_pio_s1;
  input            button_pio_s1_irq;
  input   [  2: 0] button_pio_s1_readdata;
  input            clk;
  input   [ 22: 0] pb_cpu_to_io_m1_address_to_slave;
  input            pb_cpu_to_io_m1_burstcount;
  input            pb_cpu_to_io_m1_chipselect;
  input            pb_cpu_to_io_m1_latency_counter;
  input            pb_cpu_to_io_m1_read;
  input            pb_cpu_to_io_m1_write;
  input   [ 31: 0] pb_cpu_to_io_m1_writedata;
  input            reset_n;

  wire    [  1: 0] button_pio_s1_address;
  wire             button_pio_s1_allgrants;
  wire             button_pio_s1_allow_new_arb_cycle;
  wire             button_pio_s1_any_bursting_master_saved_grant;
  wire             button_pio_s1_any_continuerequest;
  wire             button_pio_s1_arb_counter_enable;
  reg              button_pio_s1_arb_share_counter;
  wire             button_pio_s1_arb_share_counter_next_value;
  wire             button_pio_s1_arb_share_set_values;
  wire             button_pio_s1_beginbursttransfer_internal;
  wire             button_pio_s1_begins_xfer;
  wire             button_pio_s1_chipselect;
  wire             button_pio_s1_end_xfer;
  wire             button_pio_s1_firsttransfer;
  wire             button_pio_s1_grant_vector;
  wire             button_pio_s1_in_a_read_cycle;
  wire             button_pio_s1_in_a_write_cycle;
  wire             button_pio_s1_irq_from_sa;
  wire             button_pio_s1_master_qreq_vector;
  wire             button_pio_s1_non_bursting_master_requests;
  wire    [  2: 0] button_pio_s1_readdata_from_sa;
  reg              button_pio_s1_reg_firsttransfer;
  wire             button_pio_s1_reset_n;
  reg              button_pio_s1_slavearbiterlockenable;
  wire             button_pio_s1_slavearbiterlockenable2;
  wire             button_pio_s1_unreg_firsttransfer;
  wire             button_pio_s1_waits_for_read;
  wire             button_pio_s1_waits_for_write;
  wire             button_pio_s1_write_n;
  wire    [  2: 0] button_pio_s1_writedata;
  reg              d1_button_pio_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_button_pio_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             pb_cpu_to_io_m1_arbiterlock;
  wire             pb_cpu_to_io_m1_arbiterlock2;
  wire             pb_cpu_to_io_m1_continuerequest;
  wire             pb_cpu_to_io_m1_granted_button_pio_s1;
  wire             pb_cpu_to_io_m1_qualified_request_button_pio_s1;
  wire             pb_cpu_to_io_m1_read_data_valid_button_pio_s1;
  wire             pb_cpu_to_io_m1_requests_button_pio_s1;
  wire             pb_cpu_to_io_m1_saved_grant_button_pio_s1;
  wire    [ 22: 0] shifted_address_to_button_pio_s1_from_pb_cpu_to_io_m1;
  wire             wait_for_button_pio_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~button_pio_s1_end_xfer;
    end


  assign button_pio_s1_begins_xfer = ~d1_reasons_to_wait & ((pb_cpu_to_io_m1_qualified_request_button_pio_s1));
  //assign button_pio_s1_readdata_from_sa = button_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign button_pio_s1_readdata_from_sa = button_pio_s1_readdata;

  assign pb_cpu_to_io_m1_requests_button_pio_s1 = ({pb_cpu_to_io_m1_address_to_slave[22 : 4] , 4'b0} == 23'h4d00) & pb_cpu_to_io_m1_chipselect;
  //button_pio_s1_arb_share_counter set values, which is an e_mux
  assign button_pio_s1_arb_share_set_values = 1;

  //button_pio_s1_non_bursting_master_requests mux, which is an e_mux
  assign button_pio_s1_non_bursting_master_requests = pb_cpu_to_io_m1_requests_button_pio_s1;

  //button_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign button_pio_s1_any_bursting_master_saved_grant = 0;

  //button_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign button_pio_s1_arb_share_counter_next_value = button_pio_s1_firsttransfer ? (button_pio_s1_arb_share_set_values - 1) : |button_pio_s1_arb_share_counter ? (button_pio_s1_arb_share_counter - 1) : 0;

  //button_pio_s1_allgrants all slave grants, which is an e_mux
  assign button_pio_s1_allgrants = |button_pio_s1_grant_vector;

  //button_pio_s1_end_xfer assignment, which is an e_assign
  assign button_pio_s1_end_xfer = ~(button_pio_s1_waits_for_read | button_pio_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_button_pio_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_button_pio_s1 = button_pio_s1_end_xfer & (~button_pio_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //button_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign button_pio_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_button_pio_s1 & button_pio_s1_allgrants) | (end_xfer_arb_share_counter_term_button_pio_s1 & ~button_pio_s1_non_bursting_master_requests);

  //button_pio_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          button_pio_s1_arb_share_counter <= 0;
      else if (button_pio_s1_arb_counter_enable)
          button_pio_s1_arb_share_counter <= button_pio_s1_arb_share_counter_next_value;
    end


  //button_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          button_pio_s1_slavearbiterlockenable <= 0;
      else if ((|button_pio_s1_master_qreq_vector & end_xfer_arb_share_counter_term_button_pio_s1) | (end_xfer_arb_share_counter_term_button_pio_s1 & ~button_pio_s1_non_bursting_master_requests))
          button_pio_s1_slavearbiterlockenable <= |button_pio_s1_arb_share_counter_next_value;
    end


  //pb_cpu_to_io/m1 button_pio/s1 arbiterlock, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock = button_pio_s1_slavearbiterlockenable & pb_cpu_to_io_m1_continuerequest;

  //button_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign button_pio_s1_slavearbiterlockenable2 = |button_pio_s1_arb_share_counter_next_value;

  //pb_cpu_to_io/m1 button_pio/s1 arbiterlock2, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock2 = button_pio_s1_slavearbiterlockenable2 & pb_cpu_to_io_m1_continuerequest;

  //button_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign button_pio_s1_any_continuerequest = 1;

  //pb_cpu_to_io_m1_continuerequest continued request, which is an e_assign
  assign pb_cpu_to_io_m1_continuerequest = 1;

  assign pb_cpu_to_io_m1_qualified_request_button_pio_s1 = pb_cpu_to_io_m1_requests_button_pio_s1 & ~(((pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ((pb_cpu_to_io_m1_latency_counter != 0))));
  //local readdatavalid pb_cpu_to_io_m1_read_data_valid_button_pio_s1, which is an e_mux
  assign pb_cpu_to_io_m1_read_data_valid_button_pio_s1 = pb_cpu_to_io_m1_granted_button_pio_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ~button_pio_s1_waits_for_read;

  //button_pio_s1_writedata mux, which is an e_mux
  assign button_pio_s1_writedata = pb_cpu_to_io_m1_writedata;

  //master is always granted when requested
  assign pb_cpu_to_io_m1_granted_button_pio_s1 = pb_cpu_to_io_m1_qualified_request_button_pio_s1;

  //pb_cpu_to_io/m1 saved-grant button_pio/s1, which is an e_assign
  assign pb_cpu_to_io_m1_saved_grant_button_pio_s1 = pb_cpu_to_io_m1_requests_button_pio_s1;

  //allow new arb cycle for button_pio/s1, which is an e_assign
  assign button_pio_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign button_pio_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign button_pio_s1_master_qreq_vector = 1;

  //button_pio_s1_reset_n assignment, which is an e_assign
  assign button_pio_s1_reset_n = reset_n;

  assign button_pio_s1_chipselect = pb_cpu_to_io_m1_granted_button_pio_s1;
  //button_pio_s1_firsttransfer first transaction, which is an e_assign
  assign button_pio_s1_firsttransfer = button_pio_s1_begins_xfer ? button_pio_s1_unreg_firsttransfer : button_pio_s1_reg_firsttransfer;

  //button_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign button_pio_s1_unreg_firsttransfer = ~(button_pio_s1_slavearbiterlockenable & button_pio_s1_any_continuerequest);

  //button_pio_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          button_pio_s1_reg_firsttransfer <= 1'b1;
      else if (button_pio_s1_begins_xfer)
          button_pio_s1_reg_firsttransfer <= button_pio_s1_unreg_firsttransfer;
    end


  //button_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign button_pio_s1_beginbursttransfer_internal = button_pio_s1_begins_xfer;

  //~button_pio_s1_write_n assignment, which is an e_mux
  assign button_pio_s1_write_n = ~(pb_cpu_to_io_m1_granted_button_pio_s1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect));

  assign shifted_address_to_button_pio_s1_from_pb_cpu_to_io_m1 = pb_cpu_to_io_m1_address_to_slave;
  //button_pio_s1_address mux, which is an e_mux
  assign button_pio_s1_address = shifted_address_to_button_pio_s1_from_pb_cpu_to_io_m1 >> 2;

  //d1_button_pio_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_button_pio_s1_end_xfer <= 1;
      else 
        d1_button_pio_s1_end_xfer <= button_pio_s1_end_xfer;
    end


  //button_pio_s1_waits_for_read in a cycle, which is an e_mux
  assign button_pio_s1_waits_for_read = button_pio_s1_in_a_read_cycle & button_pio_s1_begins_xfer;

  //button_pio_s1_in_a_read_cycle assignment, which is an e_assign
  assign button_pio_s1_in_a_read_cycle = pb_cpu_to_io_m1_granted_button_pio_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = button_pio_s1_in_a_read_cycle;

  //button_pio_s1_waits_for_write in a cycle, which is an e_mux
  assign button_pio_s1_waits_for_write = button_pio_s1_in_a_write_cycle & 0;

  //button_pio_s1_in_a_write_cycle assignment, which is an e_assign
  assign button_pio_s1_in_a_write_cycle = pb_cpu_to_io_m1_granted_button_pio_s1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = button_pio_s1_in_a_write_cycle;

  assign wait_for_button_pio_s1_counter = 0;
  //assign button_pio_s1_irq_from_sa = button_pio_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign button_pio_s1_irq_from_sa = button_pio_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //button_pio/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pb_cpu_to_io/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_io_m1_requests_button_pio_s1 && (pb_cpu_to_io_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pb_cpu_to_io/m1 drove 0 on its 'burstcount' port while accessing slave button_pio/s1", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_jtag_debug_module_arbitrator (
                                          // inputs:
                                           clk,
                                           cpu_data_master_address_to_slave,
                                           cpu_data_master_byteenable,
                                           cpu_data_master_debugaccess,
                                           cpu_data_master_latency_counter,
                                           cpu_data_master_read,
                                           cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register,
                                           cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register,
                                           cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register,
                                           cpu_data_master_write,
                                           cpu_data_master_writedata,
                                           cpu_instruction_master_address_to_slave,
                                           cpu_instruction_master_latency_counter,
                                           cpu_instruction_master_read,
                                           cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register,
                                           cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register,
                                           cpu_jtag_debug_module_readdata,
                                           cpu_jtag_debug_module_resetrequest,
                                           reset_n,

                                          // outputs:
                                           cpu_data_master_granted_cpu_jtag_debug_module,
                                           cpu_data_master_qualified_request_cpu_jtag_debug_module,
                                           cpu_data_master_read_data_valid_cpu_jtag_debug_module,
                                           cpu_data_master_requests_cpu_jtag_debug_module,
                                           cpu_instruction_master_granted_cpu_jtag_debug_module,
                                           cpu_instruction_master_qualified_request_cpu_jtag_debug_module,
                                           cpu_instruction_master_read_data_valid_cpu_jtag_debug_module,
                                           cpu_instruction_master_requests_cpu_jtag_debug_module,
                                           cpu_jtag_debug_module_address,
                                           cpu_jtag_debug_module_begintransfer,
                                           cpu_jtag_debug_module_byteenable,
                                           cpu_jtag_debug_module_chipselect,
                                           cpu_jtag_debug_module_debugaccess,
                                           cpu_jtag_debug_module_readdata_from_sa,
                                           cpu_jtag_debug_module_reset_n,
                                           cpu_jtag_debug_module_resetrequest_from_sa,
                                           cpu_jtag_debug_module_write,
                                           cpu_jtag_debug_module_writedata,
                                           d1_cpu_jtag_debug_module_end_xfer
                                        )
;

  output           cpu_data_master_granted_cpu_jtag_debug_module;
  output           cpu_data_master_qualified_request_cpu_jtag_debug_module;
  output           cpu_data_master_read_data_valid_cpu_jtag_debug_module;
  output           cpu_data_master_requests_cpu_jtag_debug_module;
  output           cpu_instruction_master_granted_cpu_jtag_debug_module;
  output           cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  output           cpu_instruction_master_read_data_valid_cpu_jtag_debug_module;
  output           cpu_instruction_master_requests_cpu_jtag_debug_module;
  output  [  8: 0] cpu_jtag_debug_module_address;
  output           cpu_jtag_debug_module_begintransfer;
  output  [  3: 0] cpu_jtag_debug_module_byteenable;
  output           cpu_jtag_debug_module_chipselect;
  output           cpu_jtag_debug_module_debugaccess;
  output  [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  output           cpu_jtag_debug_module_reset_n;
  output           cpu_jtag_debug_module_resetrequest_from_sa;
  output           cpu_jtag_debug_module_write;
  output  [ 31: 0] cpu_jtag_debug_module_writedata;
  output           d1_cpu_jtag_debug_module_end_xfer;
  input            clk;
  input   [ 28: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register;
  input            cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register;
  input            cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 28: 0] cpu_instruction_master_address_to_slave;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register;
  input            cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register;
  input   [ 31: 0] cpu_jtag_debug_module_readdata;
  input            cpu_jtag_debug_module_resetrequest;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_cpu_jtag_debug_module;
  wire             cpu_data_master_qualified_request_cpu_jtag_debug_module;
  wire             cpu_data_master_read_data_valid_cpu_jtag_debug_module;
  wire             cpu_data_master_requests_cpu_jtag_debug_module;
  wire             cpu_data_master_saved_grant_cpu_jtag_debug_module;
  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_cpu_jtag_debug_module;
  wire             cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  wire             cpu_instruction_master_read_data_valid_cpu_jtag_debug_module;
  wire             cpu_instruction_master_requests_cpu_jtag_debug_module;
  wire             cpu_instruction_master_saved_grant_cpu_jtag_debug_module;
  wire    [  8: 0] cpu_jtag_debug_module_address;
  wire             cpu_jtag_debug_module_allgrants;
  wire             cpu_jtag_debug_module_allow_new_arb_cycle;
  wire             cpu_jtag_debug_module_any_bursting_master_saved_grant;
  wire             cpu_jtag_debug_module_any_continuerequest;
  reg     [  1: 0] cpu_jtag_debug_module_arb_addend;
  wire             cpu_jtag_debug_module_arb_counter_enable;
  reg              cpu_jtag_debug_module_arb_share_counter;
  wire             cpu_jtag_debug_module_arb_share_counter_next_value;
  wire             cpu_jtag_debug_module_arb_share_set_values;
  wire    [  1: 0] cpu_jtag_debug_module_arb_winner;
  wire             cpu_jtag_debug_module_arbitration_holdoff_internal;
  wire             cpu_jtag_debug_module_beginbursttransfer_internal;
  wire             cpu_jtag_debug_module_begins_xfer;
  wire             cpu_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_jtag_debug_module_byteenable;
  wire             cpu_jtag_debug_module_chipselect;
  wire    [  3: 0] cpu_jtag_debug_module_chosen_master_double_vector;
  wire    [  1: 0] cpu_jtag_debug_module_chosen_master_rot_left;
  wire             cpu_jtag_debug_module_debugaccess;
  wire             cpu_jtag_debug_module_end_xfer;
  wire             cpu_jtag_debug_module_firsttransfer;
  wire    [  1: 0] cpu_jtag_debug_module_grant_vector;
  wire             cpu_jtag_debug_module_in_a_read_cycle;
  wire             cpu_jtag_debug_module_in_a_write_cycle;
  wire    [  1: 0] cpu_jtag_debug_module_master_qreq_vector;
  wire             cpu_jtag_debug_module_non_bursting_master_requests;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  reg              cpu_jtag_debug_module_reg_firsttransfer;
  wire             cpu_jtag_debug_module_reset_n;
  wire             cpu_jtag_debug_module_resetrequest_from_sa;
  reg     [  1: 0] cpu_jtag_debug_module_saved_chosen_master_vector;
  reg              cpu_jtag_debug_module_slavearbiterlockenable;
  wire             cpu_jtag_debug_module_slavearbiterlockenable2;
  wire             cpu_jtag_debug_module_unreg_firsttransfer;
  wire             cpu_jtag_debug_module_waits_for_read;
  wire             cpu_jtag_debug_module_waits_for_write;
  wire             cpu_jtag_debug_module_write;
  wire    [ 31: 0] cpu_jtag_debug_module_writedata;
  reg              d1_cpu_jtag_debug_module_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_cpu_jtag_debug_module;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module;
  reg              last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module;
  wire    [ 28: 0] shifted_address_to_cpu_jtag_debug_module_from_cpu_data_master;
  wire    [ 28: 0] shifted_address_to_cpu_jtag_debug_module_from_cpu_instruction_master;
  wire             wait_for_cpu_jtag_debug_module_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~cpu_jtag_debug_module_end_xfer;
    end


  assign cpu_jtag_debug_module_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_cpu_jtag_debug_module | cpu_instruction_master_qualified_request_cpu_jtag_debug_module));
  //assign cpu_jtag_debug_module_readdata_from_sa = cpu_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_jtag_debug_module_readdata_from_sa = cpu_jtag_debug_module_readdata;

  assign cpu_data_master_requests_cpu_jtag_debug_module = ({cpu_data_master_address_to_slave[28 : 11] , 11'b0} == 29'h7fff800) & (cpu_data_master_read | cpu_data_master_write);
  //cpu_jtag_debug_module_arb_share_counter set values, which is an e_mux
  assign cpu_jtag_debug_module_arb_share_set_values = 1;

  //cpu_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  assign cpu_jtag_debug_module_non_bursting_master_requests = cpu_data_master_requests_cpu_jtag_debug_module |
    cpu_instruction_master_requests_cpu_jtag_debug_module |
    cpu_data_master_requests_cpu_jtag_debug_module |
    cpu_instruction_master_requests_cpu_jtag_debug_module;

  //cpu_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  assign cpu_jtag_debug_module_any_bursting_master_saved_grant = 0;

  //cpu_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  assign cpu_jtag_debug_module_arb_share_counter_next_value = cpu_jtag_debug_module_firsttransfer ? (cpu_jtag_debug_module_arb_share_set_values - 1) : |cpu_jtag_debug_module_arb_share_counter ? (cpu_jtag_debug_module_arb_share_counter - 1) : 0;

  //cpu_jtag_debug_module_allgrants all slave grants, which is an e_mux
  assign cpu_jtag_debug_module_allgrants = (|cpu_jtag_debug_module_grant_vector) |
    (|cpu_jtag_debug_module_grant_vector) |
    (|cpu_jtag_debug_module_grant_vector) |
    (|cpu_jtag_debug_module_grant_vector);

  //cpu_jtag_debug_module_end_xfer assignment, which is an e_assign
  assign cpu_jtag_debug_module_end_xfer = ~(cpu_jtag_debug_module_waits_for_read | cpu_jtag_debug_module_waits_for_write);

  //end_xfer_arb_share_counter_term_cpu_jtag_debug_module arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_cpu_jtag_debug_module = cpu_jtag_debug_module_end_xfer & (~cpu_jtag_debug_module_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //cpu_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  assign cpu_jtag_debug_module_arb_counter_enable = (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & cpu_jtag_debug_module_allgrants) | (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & ~cpu_jtag_debug_module_non_bursting_master_requests);

  //cpu_jtag_debug_module_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_arb_share_counter <= 0;
      else if (cpu_jtag_debug_module_arb_counter_enable)
          cpu_jtag_debug_module_arb_share_counter <= cpu_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_slavearbiterlockenable <= 0;
      else if ((|cpu_jtag_debug_module_master_qreq_vector & end_xfer_arb_share_counter_term_cpu_jtag_debug_module) | (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & ~cpu_jtag_debug_module_non_bursting_master_requests))
          cpu_jtag_debug_module_slavearbiterlockenable <= |cpu_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu/data_master cpu/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = cpu_jtag_debug_module_slavearbiterlockenable & cpu_data_master_continuerequest;

  //cpu_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign cpu_jtag_debug_module_slavearbiterlockenable2 = |cpu_jtag_debug_module_arb_share_counter_next_value;

  //cpu/data_master cpu/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = cpu_jtag_debug_module_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //cpu/instruction_master cpu/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = cpu_jtag_debug_module_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //cpu/instruction_master cpu/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = cpu_jtag_debug_module_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //cpu/instruction_master granted cpu/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module <= cpu_instruction_master_saved_grant_cpu_jtag_debug_module ? 1 : (cpu_jtag_debug_module_arbitration_holdoff_internal | ~cpu_instruction_master_requests_cpu_jtag_debug_module) ? 0 : last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module;
    end


  //cpu_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_instruction_master_continuerequest = last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module & cpu_instruction_master_requests_cpu_jtag_debug_module;

  //cpu_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  assign cpu_jtag_debug_module_any_continuerequest = cpu_instruction_master_continuerequest |
    cpu_data_master_continuerequest;

  assign cpu_data_master_qualified_request_cpu_jtag_debug_module = cpu_data_master_requests_cpu_jtag_debug_module & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (|cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register) | (|cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register) | (|cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register))) | cpu_instruction_master_arbiterlock);
  //local readdatavalid cpu_data_master_read_data_valid_cpu_jtag_debug_module, which is an e_mux
  assign cpu_data_master_read_data_valid_cpu_jtag_debug_module = cpu_data_master_granted_cpu_jtag_debug_module & cpu_data_master_read & ~cpu_jtag_debug_module_waits_for_read;

  //cpu_jtag_debug_module_writedata mux, which is an e_mux
  assign cpu_jtag_debug_module_writedata = cpu_data_master_writedata;

  assign cpu_instruction_master_requests_cpu_jtag_debug_module = (({cpu_instruction_master_address_to_slave[28 : 11] , 11'b0} == 29'h7fff800) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //cpu/data_master granted cpu/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module <= cpu_data_master_saved_grant_cpu_jtag_debug_module ? 1 : (cpu_jtag_debug_module_arbitration_holdoff_internal | ~cpu_data_master_requests_cpu_jtag_debug_module) ? 0 : last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module;
    end


  //cpu_data_master_continuerequest continued request, which is an e_mux
  assign cpu_data_master_continuerequest = last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module & cpu_data_master_requests_cpu_jtag_debug_module;

  assign cpu_instruction_master_qualified_request_cpu_jtag_debug_module = cpu_instruction_master_requests_cpu_jtag_debug_module & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (|cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register) | (|cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register))) | cpu_data_master_arbiterlock);
  //local readdatavalid cpu_instruction_master_read_data_valid_cpu_jtag_debug_module, which is an e_mux
  assign cpu_instruction_master_read_data_valid_cpu_jtag_debug_module = cpu_instruction_master_granted_cpu_jtag_debug_module & cpu_instruction_master_read & ~cpu_jtag_debug_module_waits_for_read;

  //allow new arb cycle for cpu/jtag_debug_module, which is an e_assign
  assign cpu_jtag_debug_module_allow_new_arb_cycle = ~cpu_data_master_arbiterlock & ~cpu_instruction_master_arbiterlock;

  //cpu/instruction_master assignment into master qualified-requests vector for cpu/jtag_debug_module, which is an e_assign
  assign cpu_jtag_debug_module_master_qreq_vector[0] = cpu_instruction_master_qualified_request_cpu_jtag_debug_module;

  //cpu/instruction_master grant cpu/jtag_debug_module, which is an e_assign
  assign cpu_instruction_master_granted_cpu_jtag_debug_module = cpu_jtag_debug_module_grant_vector[0];

  //cpu/instruction_master saved-grant cpu/jtag_debug_module, which is an e_assign
  assign cpu_instruction_master_saved_grant_cpu_jtag_debug_module = cpu_jtag_debug_module_arb_winner[0] && cpu_instruction_master_requests_cpu_jtag_debug_module;

  //cpu/data_master assignment into master qualified-requests vector for cpu/jtag_debug_module, which is an e_assign
  assign cpu_jtag_debug_module_master_qreq_vector[1] = cpu_data_master_qualified_request_cpu_jtag_debug_module;

  //cpu/data_master grant cpu/jtag_debug_module, which is an e_assign
  assign cpu_data_master_granted_cpu_jtag_debug_module = cpu_jtag_debug_module_grant_vector[1];

  //cpu/data_master saved-grant cpu/jtag_debug_module, which is an e_assign
  assign cpu_data_master_saved_grant_cpu_jtag_debug_module = cpu_jtag_debug_module_arb_winner[1] && cpu_data_master_requests_cpu_jtag_debug_module;

  //cpu/jtag_debug_module chosen-master double-vector, which is an e_assign
  assign cpu_jtag_debug_module_chosen_master_double_vector = {cpu_jtag_debug_module_master_qreq_vector, cpu_jtag_debug_module_master_qreq_vector} & ({~cpu_jtag_debug_module_master_qreq_vector, ~cpu_jtag_debug_module_master_qreq_vector} + cpu_jtag_debug_module_arb_addend);

  //stable onehot encoding of arb winner
  assign cpu_jtag_debug_module_arb_winner = (cpu_jtag_debug_module_allow_new_arb_cycle & | cpu_jtag_debug_module_grant_vector) ? cpu_jtag_debug_module_grant_vector : cpu_jtag_debug_module_saved_chosen_master_vector;

  //saved cpu_jtag_debug_module_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_saved_chosen_master_vector <= 0;
      else if (cpu_jtag_debug_module_allow_new_arb_cycle)
          cpu_jtag_debug_module_saved_chosen_master_vector <= |cpu_jtag_debug_module_grant_vector ? cpu_jtag_debug_module_grant_vector : cpu_jtag_debug_module_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign cpu_jtag_debug_module_grant_vector = {(cpu_jtag_debug_module_chosen_master_double_vector[1] | cpu_jtag_debug_module_chosen_master_double_vector[3]),
    (cpu_jtag_debug_module_chosen_master_double_vector[0] | cpu_jtag_debug_module_chosen_master_double_vector[2])};

  //cpu/jtag_debug_module chosen master rotated left, which is an e_assign
  assign cpu_jtag_debug_module_chosen_master_rot_left = (cpu_jtag_debug_module_arb_winner << 1) ? (cpu_jtag_debug_module_arb_winner << 1) : 1;

  //cpu/jtag_debug_module's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_arb_addend <= 1;
      else if (|cpu_jtag_debug_module_grant_vector)
          cpu_jtag_debug_module_arb_addend <= cpu_jtag_debug_module_end_xfer? cpu_jtag_debug_module_chosen_master_rot_left : cpu_jtag_debug_module_grant_vector;
    end


  assign cpu_jtag_debug_module_begintransfer = cpu_jtag_debug_module_begins_xfer;
  //cpu_jtag_debug_module_reset_n assignment, which is an e_assign
  assign cpu_jtag_debug_module_reset_n = reset_n;

  //assign cpu_jtag_debug_module_resetrequest_from_sa = cpu_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_jtag_debug_module_resetrequest_from_sa = cpu_jtag_debug_module_resetrequest;

  assign cpu_jtag_debug_module_chipselect = cpu_data_master_granted_cpu_jtag_debug_module | cpu_instruction_master_granted_cpu_jtag_debug_module;
  //cpu_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  assign cpu_jtag_debug_module_firsttransfer = cpu_jtag_debug_module_begins_xfer ? cpu_jtag_debug_module_unreg_firsttransfer : cpu_jtag_debug_module_reg_firsttransfer;

  //cpu_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  assign cpu_jtag_debug_module_unreg_firsttransfer = ~(cpu_jtag_debug_module_slavearbiterlockenable & cpu_jtag_debug_module_any_continuerequest);

  //cpu_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_reg_firsttransfer <= 1'b1;
      else if (cpu_jtag_debug_module_begins_xfer)
          cpu_jtag_debug_module_reg_firsttransfer <= cpu_jtag_debug_module_unreg_firsttransfer;
    end


  //cpu_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign cpu_jtag_debug_module_beginbursttransfer_internal = cpu_jtag_debug_module_begins_xfer;

  //cpu_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign cpu_jtag_debug_module_arbitration_holdoff_internal = cpu_jtag_debug_module_begins_xfer & cpu_jtag_debug_module_firsttransfer;

  //cpu_jtag_debug_module_write assignment, which is an e_mux
  assign cpu_jtag_debug_module_write = cpu_data_master_granted_cpu_jtag_debug_module & cpu_data_master_write;

  assign shifted_address_to_cpu_jtag_debug_module_from_cpu_data_master = cpu_data_master_address_to_slave;
  //cpu_jtag_debug_module_address mux, which is an e_mux
  assign cpu_jtag_debug_module_address = (cpu_data_master_granted_cpu_jtag_debug_module)? (shifted_address_to_cpu_jtag_debug_module_from_cpu_data_master >> 2) :
    (shifted_address_to_cpu_jtag_debug_module_from_cpu_instruction_master >> 2);

  assign shifted_address_to_cpu_jtag_debug_module_from_cpu_instruction_master = cpu_instruction_master_address_to_slave;
  //d1_cpu_jtag_debug_module_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_cpu_jtag_debug_module_end_xfer <= 1;
      else 
        d1_cpu_jtag_debug_module_end_xfer <= cpu_jtag_debug_module_end_xfer;
    end


  //cpu_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  assign cpu_jtag_debug_module_waits_for_read = cpu_jtag_debug_module_in_a_read_cycle & cpu_jtag_debug_module_begins_xfer;

  //cpu_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  assign cpu_jtag_debug_module_in_a_read_cycle = (cpu_data_master_granted_cpu_jtag_debug_module & cpu_data_master_read) | (cpu_instruction_master_granted_cpu_jtag_debug_module & cpu_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cpu_jtag_debug_module_in_a_read_cycle;

  //cpu_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  assign cpu_jtag_debug_module_waits_for_write = cpu_jtag_debug_module_in_a_write_cycle & 0;

  //cpu_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  assign cpu_jtag_debug_module_in_a_write_cycle = cpu_data_master_granted_cpu_jtag_debug_module & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cpu_jtag_debug_module_in_a_write_cycle;

  assign wait_for_cpu_jtag_debug_module_counter = 0;
  //cpu_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  assign cpu_jtag_debug_module_byteenable = (cpu_data_master_granted_cpu_jtag_debug_module)? cpu_data_master_byteenable :
    -1;

  //debugaccess mux, which is an e_mux
  assign cpu_jtag_debug_module_debugaccess = (cpu_data_master_granted_cpu_jtag_debug_module)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu/jtag_debug_module enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_granted_cpu_jtag_debug_module + cpu_instruction_master_granted_cpu_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_saved_grant_cpu_jtag_debug_module + cpu_instruction_master_saved_grant_cpu_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_data_master_arbitrator (
                                    // inputs:
                                     button_pio_s1_irq_from_sa,
                                     clk,
                                     cpu_data_master_address,
                                     cpu_data_master_byteenable,
                                     cpu_data_master_granted_cpu_jtag_debug_module,
                                     cpu_data_master_granted_pb_cpu_to_ddr3_top_s1,
                                     cpu_data_master_granted_pb_cpu_to_fsm_s1,
                                     cpu_data_master_granted_pb_cpu_to_io_s1,
                                     cpu_data_master_qualified_request_cpu_jtag_debug_module,
                                     cpu_data_master_qualified_request_pb_cpu_to_ddr3_top_s1,
                                     cpu_data_master_qualified_request_pb_cpu_to_fsm_s1,
                                     cpu_data_master_qualified_request_pb_cpu_to_io_s1,
                                     cpu_data_master_read,
                                     cpu_data_master_read_data_valid_cpu_jtag_debug_module,
                                     cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1,
                                     cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register,
                                     cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1,
                                     cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register,
                                     cpu_data_master_read_data_valid_pb_cpu_to_io_s1,
                                     cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register,
                                     cpu_data_master_requests_cpu_jtag_debug_module,
                                     cpu_data_master_requests_pb_cpu_to_ddr3_top_s1,
                                     cpu_data_master_requests_pb_cpu_to_fsm_s1,
                                     cpu_data_master_requests_pb_cpu_to_io_s1,
                                     cpu_data_master_write,
                                     cpu_data_master_writedata,
                                     cpu_jtag_debug_module_readdata_from_sa,
                                     d1_cpu_jtag_debug_module_end_xfer,
                                     d1_pb_cpu_to_ddr3_top_s1_end_xfer,
                                     d1_pb_cpu_to_fsm_s1_end_xfer,
                                     d1_pb_cpu_to_io_s1_end_xfer,
                                     dipsw_pio_s1_irq_from_sa,
                                     jtag_uart_avalon_jtag_slave_irq_from_sa,
                                     pb_cpu_to_ddr3_top_s1_readdata_from_sa,
                                     pb_cpu_to_ddr3_top_s1_waitrequest_from_sa,
                                     pb_cpu_to_fsm_s1_readdata_from_sa,
                                     pb_cpu_to_fsm_s1_waitrequest_from_sa,
                                     pb_cpu_to_io_s1_readdata_from_sa,
                                     pb_cpu_to_io_s1_waitrequest_from_sa,
                                     reset_n,
                                     sgdma_rx_csr_irq_from_sa,
                                     sgdma_tx_csr_irq_from_sa,
                                     timer_1ms_s1_irq_from_sa,
                                     uart_s1_irq_from_sa,

                                    // outputs:
                                     cpu_data_master_address_to_slave,
                                     cpu_data_master_irq,
                                     cpu_data_master_latency_counter,
                                     cpu_data_master_readdata,
                                     cpu_data_master_readdatavalid,
                                     cpu_data_master_waitrequest
                                  )
;

  output  [ 28: 0] cpu_data_master_address_to_slave;
  output  [ 31: 0] cpu_data_master_irq;
  output           cpu_data_master_latency_counter;
  output  [ 31: 0] cpu_data_master_readdata;
  output           cpu_data_master_readdatavalid;
  output           cpu_data_master_waitrequest;
  input            button_pio_s1_irq_from_sa;
  input            clk;
  input   [ 28: 0] cpu_data_master_address;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_granted_cpu_jtag_debug_module;
  input            cpu_data_master_granted_pb_cpu_to_ddr3_top_s1;
  input            cpu_data_master_granted_pb_cpu_to_fsm_s1;
  input            cpu_data_master_granted_pb_cpu_to_io_s1;
  input            cpu_data_master_qualified_request_cpu_jtag_debug_module;
  input            cpu_data_master_qualified_request_pb_cpu_to_ddr3_top_s1;
  input            cpu_data_master_qualified_request_pb_cpu_to_fsm_s1;
  input            cpu_data_master_qualified_request_pb_cpu_to_io_s1;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_cpu_jtag_debug_module;
  input            cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1;
  input            cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register;
  input            cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1;
  input            cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register;
  input            cpu_data_master_read_data_valid_pb_cpu_to_io_s1;
  input            cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register;
  input            cpu_data_master_requests_cpu_jtag_debug_module;
  input            cpu_data_master_requests_pb_cpu_to_ddr3_top_s1;
  input            cpu_data_master_requests_pb_cpu_to_fsm_s1;
  input            cpu_data_master_requests_pb_cpu_to_io_s1;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_jtag_debug_module_end_xfer;
  input            d1_pb_cpu_to_ddr3_top_s1_end_xfer;
  input            d1_pb_cpu_to_fsm_s1_end_xfer;
  input            d1_pb_cpu_to_io_s1_end_xfer;
  input            dipsw_pio_s1_irq_from_sa;
  input            jtag_uart_avalon_jtag_slave_irq_from_sa;
  input   [ 31: 0] pb_cpu_to_ddr3_top_s1_readdata_from_sa;
  input            pb_cpu_to_ddr3_top_s1_waitrequest_from_sa;
  input   [ 31: 0] pb_cpu_to_fsm_s1_readdata_from_sa;
  input            pb_cpu_to_fsm_s1_waitrequest_from_sa;
  input   [ 31: 0] pb_cpu_to_io_s1_readdata_from_sa;
  input            pb_cpu_to_io_s1_waitrequest_from_sa;
  input            reset_n;
  input            sgdma_rx_csr_irq_from_sa;
  input            sgdma_tx_csr_irq_from_sa;
  input            timer_1ms_s1_irq_from_sa;
  input            uart_s1_irq_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 28: 0] cpu_data_master_address_last_time;
  wire    [ 28: 0] cpu_data_master_address_to_slave;
  reg     [  3: 0] cpu_data_master_byteenable_last_time;
  wire    [ 31: 0] cpu_data_master_irq;
  wire             cpu_data_master_is_granted_some_slave;
  reg              cpu_data_master_latency_counter;
  reg              cpu_data_master_read_but_no_slave_selected;
  reg              cpu_data_master_read_last_time;
  wire    [ 31: 0] cpu_data_master_readdata;
  wire             cpu_data_master_readdatavalid;
  wire             cpu_data_master_run;
  wire             cpu_data_master_waitrequest;
  reg              cpu_data_master_write_last_time;
  reg     [ 31: 0] cpu_data_master_writedata_last_time;
  wire             latency_load_value;
  wire             p1_cpu_data_master_latency_counter;
  wire             pre_flush_cpu_data_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_data_master_qualified_request_cpu_jtag_debug_module | ~cpu_data_master_requests_cpu_jtag_debug_module) & (cpu_data_master_granted_cpu_jtag_debug_module | ~cpu_data_master_qualified_request_cpu_jtag_debug_module) & ((~cpu_data_master_qualified_request_cpu_jtag_debug_module | ~cpu_data_master_read | (1 & ~d1_cpu_jtag_debug_module_end_xfer & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_cpu_jtag_debug_module | ~cpu_data_master_write | (1 & cpu_data_master_write)));

  //cascaded wait assignment, which is an e_assign
  assign cpu_data_master_run = r_0 & r_1;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_data_master_qualified_request_pb_cpu_to_ddr3_top_s1 | ~cpu_data_master_requests_pb_cpu_to_ddr3_top_s1) & (cpu_data_master_granted_pb_cpu_to_ddr3_top_s1 | ~cpu_data_master_qualified_request_pb_cpu_to_ddr3_top_s1) & ((~cpu_data_master_qualified_request_pb_cpu_to_ddr3_top_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~pb_cpu_to_ddr3_top_s1_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_pb_cpu_to_ddr3_top_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~pb_cpu_to_ddr3_top_s1_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_pb_cpu_to_fsm_s1 | ~cpu_data_master_requests_pb_cpu_to_fsm_s1) & (cpu_data_master_granted_pb_cpu_to_fsm_s1 | ~cpu_data_master_qualified_request_pb_cpu_to_fsm_s1) & ((~cpu_data_master_qualified_request_pb_cpu_to_fsm_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~pb_cpu_to_fsm_s1_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_pb_cpu_to_fsm_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~pb_cpu_to_fsm_s1_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_pb_cpu_to_io_s1 | ~cpu_data_master_requests_pb_cpu_to_io_s1) & ((~cpu_data_master_qualified_request_pb_cpu_to_io_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~pb_cpu_to_io_s1_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_pb_cpu_to_io_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~pb_cpu_to_io_s1_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write))));

  //irq assign, which is an e_assign
  assign cpu_data_master_irq = {1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    timer_1ms_s1_irq_from_sa,
    uart_s1_irq_from_sa,
    button_pio_s1_irq_from_sa,
    dipsw_pio_s1_irq_from_sa,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    sgdma_tx_csr_irq_from_sa,
    sgdma_rx_csr_irq_from_sa,
    jtag_uart_avalon_jtag_slave_irq_from_sa,
    1'b0};

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_data_master_address_to_slave = cpu_data_master_address[28 : 0];

  //cpu_data_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_read_but_no_slave_selected <= 0;
      else 
        cpu_data_master_read_but_no_slave_selected <= cpu_data_master_read & cpu_data_master_run & ~cpu_data_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_data_master_is_granted_some_slave = cpu_data_master_granted_cpu_jtag_debug_module |
    cpu_data_master_granted_pb_cpu_to_ddr3_top_s1 |
    cpu_data_master_granted_pb_cpu_to_fsm_s1 |
    cpu_data_master_granted_pb_cpu_to_io_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_data_master_readdatavalid = cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1 |
    cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1 |
    cpu_data_master_read_data_valid_pb_cpu_to_io_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_data_master_readdatavalid = cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_data_valid_cpu_jtag_debug_module |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid;

  //cpu/data_master readdata mux, which is an e_mux
  assign cpu_data_master_readdata = ({32 {~(cpu_data_master_qualified_request_cpu_jtag_debug_module & cpu_data_master_read)}} | cpu_jtag_debug_module_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1}} | pb_cpu_to_ddr3_top_s1_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1}} | pb_cpu_to_fsm_s1_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_pb_cpu_to_io_s1}} | pb_cpu_to_io_s1_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_data_master_waitrequest = ~cpu_data_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_latency_counter <= 0;
      else 
        cpu_data_master_latency_counter <= p1_cpu_data_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_data_master_latency_counter = ((cpu_data_master_run & cpu_data_master_read))? latency_load_value :
    (cpu_data_master_latency_counter)? cpu_data_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_data_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_address_last_time <= 0;
      else 
        cpu_data_master_address_last_time <= cpu_data_master_address;
    end


  //cpu/data_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_data_master_waitrequest & (cpu_data_master_read | cpu_data_master_write);
    end


  //cpu_data_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_address != cpu_data_master_address_last_time))
        begin
          $write("%0d ns: cpu_data_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_byteenable_last_time <= 0;
      else 
        cpu_data_master_byteenable_last_time <= cpu_data_master_byteenable;
    end


  //cpu_data_master_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_byteenable != cpu_data_master_byteenable_last_time))
        begin
          $write("%0d ns: cpu_data_master_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_read_last_time <= 0;
      else 
        cpu_data_master_read_last_time <= cpu_data_master_read;
    end


  //cpu_data_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_read != cpu_data_master_read_last_time))
        begin
          $write("%0d ns: cpu_data_master_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_write_last_time <= 0;
      else 
        cpu_data_master_write_last_time <= cpu_data_master_write;
    end


  //cpu_data_master_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_write != cpu_data_master_write_last_time))
        begin
          $write("%0d ns: cpu_data_master_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_writedata_last_time <= 0;
      else 
        cpu_data_master_writedata_last_time <= cpu_data_master_writedata;
    end


  //cpu_data_master_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_writedata != cpu_data_master_writedata_last_time) & cpu_data_master_write)
        begin
          $write("%0d ns: cpu_data_master_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_instruction_master_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_instruction_master_address,
                                            cpu_instruction_master_granted_cpu_jtag_debug_module,
                                            cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1,
                                            cpu_instruction_master_granted_pb_cpu_to_fsm_s1,
                                            cpu_instruction_master_qualified_request_cpu_jtag_debug_module,
                                            cpu_instruction_master_qualified_request_pb_cpu_to_ddr3_top_s1,
                                            cpu_instruction_master_qualified_request_pb_cpu_to_fsm_s1,
                                            cpu_instruction_master_read,
                                            cpu_instruction_master_read_data_valid_cpu_jtag_debug_module,
                                            cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1,
                                            cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register,
                                            cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1,
                                            cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register,
                                            cpu_instruction_master_requests_cpu_jtag_debug_module,
                                            cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1,
                                            cpu_instruction_master_requests_pb_cpu_to_fsm_s1,
                                            cpu_jtag_debug_module_readdata_from_sa,
                                            d1_cpu_jtag_debug_module_end_xfer,
                                            d1_pb_cpu_to_ddr3_top_s1_end_xfer,
                                            d1_pb_cpu_to_fsm_s1_end_xfer,
                                            pb_cpu_to_ddr3_top_s1_readdata_from_sa,
                                            pb_cpu_to_ddr3_top_s1_waitrequest_from_sa,
                                            pb_cpu_to_fsm_s1_readdata_from_sa,
                                            pb_cpu_to_fsm_s1_waitrequest_from_sa,
                                            reset_n,

                                           // outputs:
                                            cpu_instruction_master_address_to_slave,
                                            cpu_instruction_master_latency_counter,
                                            cpu_instruction_master_readdata,
                                            cpu_instruction_master_readdatavalid,
                                            cpu_instruction_master_waitrequest
                                         )
;

  output  [ 28: 0] cpu_instruction_master_address_to_slave;
  output           cpu_instruction_master_latency_counter;
  output  [ 31: 0] cpu_instruction_master_readdata;
  output           cpu_instruction_master_readdatavalid;
  output           cpu_instruction_master_waitrequest;
  input            clk;
  input   [ 28: 0] cpu_instruction_master_address;
  input            cpu_instruction_master_granted_cpu_jtag_debug_module;
  input            cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1;
  input            cpu_instruction_master_granted_pb_cpu_to_fsm_s1;
  input            cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  input            cpu_instruction_master_qualified_request_pb_cpu_to_ddr3_top_s1;
  input            cpu_instruction_master_qualified_request_pb_cpu_to_fsm_s1;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_cpu_jtag_debug_module;
  input            cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1;
  input            cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register;
  input            cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1;
  input            cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register;
  input            cpu_instruction_master_requests_cpu_jtag_debug_module;
  input            cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1;
  input            cpu_instruction_master_requests_pb_cpu_to_fsm_s1;
  input   [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_jtag_debug_module_end_xfer;
  input            d1_pb_cpu_to_ddr3_top_s1_end_xfer;
  input            d1_pb_cpu_to_fsm_s1_end_xfer;
  input   [ 31: 0] pb_cpu_to_ddr3_top_s1_readdata_from_sa;
  input            pb_cpu_to_ddr3_top_s1_waitrequest_from_sa;
  input   [ 31: 0] pb_cpu_to_fsm_s1_readdata_from_sa;
  input            pb_cpu_to_fsm_s1_waitrequest_from_sa;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 28: 0] cpu_instruction_master_address_last_time;
  wire    [ 28: 0] cpu_instruction_master_address_to_slave;
  wire             cpu_instruction_master_is_granted_some_slave;
  reg              cpu_instruction_master_latency_counter;
  reg              cpu_instruction_master_read_but_no_slave_selected;
  reg              cpu_instruction_master_read_last_time;
  wire    [ 31: 0] cpu_instruction_master_readdata;
  wire             cpu_instruction_master_readdatavalid;
  wire             cpu_instruction_master_run;
  wire             cpu_instruction_master_waitrequest;
  wire             latency_load_value;
  wire             p1_cpu_instruction_master_latency_counter;
  wire             pre_flush_cpu_instruction_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_instruction_master_qualified_request_cpu_jtag_debug_module | ~cpu_instruction_master_requests_cpu_jtag_debug_module) & (cpu_instruction_master_granted_cpu_jtag_debug_module | ~cpu_instruction_master_qualified_request_cpu_jtag_debug_module) & ((~cpu_instruction_master_qualified_request_cpu_jtag_debug_module | ~cpu_instruction_master_read | (1 & ~d1_cpu_jtag_debug_module_end_xfer & cpu_instruction_master_read)));

  //cascaded wait assignment, which is an e_assign
  assign cpu_instruction_master_run = r_0 & r_1;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_instruction_master_qualified_request_pb_cpu_to_ddr3_top_s1 | ~cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1) & (cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1 | ~cpu_instruction_master_qualified_request_pb_cpu_to_ddr3_top_s1) & ((~cpu_instruction_master_qualified_request_pb_cpu_to_ddr3_top_s1 | ~(cpu_instruction_master_read) | (1 & ~pb_cpu_to_ddr3_top_s1_waitrequest_from_sa & (cpu_instruction_master_read)))) & 1 & (cpu_instruction_master_qualified_request_pb_cpu_to_fsm_s1 | ~cpu_instruction_master_requests_pb_cpu_to_fsm_s1) & (cpu_instruction_master_granted_pb_cpu_to_fsm_s1 | ~cpu_instruction_master_qualified_request_pb_cpu_to_fsm_s1) & ((~cpu_instruction_master_qualified_request_pb_cpu_to_fsm_s1 | ~(cpu_instruction_master_read) | (1 & ~pb_cpu_to_fsm_s1_waitrequest_from_sa & (cpu_instruction_master_read))));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_instruction_master_address_to_slave = {cpu_instruction_master_address[28],
    1'b0,
    cpu_instruction_master_address[26 : 0]};

  //cpu_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_read_but_no_slave_selected <= 0;
      else 
        cpu_instruction_master_read_but_no_slave_selected <= cpu_instruction_master_read & cpu_instruction_master_run & ~cpu_instruction_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_instruction_master_is_granted_some_slave = cpu_instruction_master_granted_cpu_jtag_debug_module |
    cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1 |
    cpu_instruction_master_granted_pb_cpu_to_fsm_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_instruction_master_readdatavalid = cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1 |
    cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_instruction_master_readdatavalid = cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid |
    cpu_instruction_master_read_data_valid_cpu_jtag_debug_module |
    cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid |
    cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid;

  //cpu/instruction_master readdata mux, which is an e_mux
  assign cpu_instruction_master_readdata = ({32 {~(cpu_instruction_master_qualified_request_cpu_jtag_debug_module & cpu_instruction_master_read)}} | cpu_jtag_debug_module_readdata_from_sa) &
    ({32 {~cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1}} | pb_cpu_to_ddr3_top_s1_readdata_from_sa) &
    ({32 {~cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1}} | pb_cpu_to_fsm_s1_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_instruction_master_waitrequest = ~cpu_instruction_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_latency_counter <= 0;
      else 
        cpu_instruction_master_latency_counter <= p1_cpu_instruction_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_instruction_master_latency_counter = ((cpu_instruction_master_run & cpu_instruction_master_read))? latency_load_value :
    (cpu_instruction_master_latency_counter)? cpu_instruction_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_instruction_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_address_last_time <= 0;
      else 
        cpu_instruction_master_address_last_time <= cpu_instruction_master_address;
    end


  //cpu/instruction_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_instruction_master_waitrequest & (cpu_instruction_master_read);
    end


  //cpu_instruction_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_instruction_master_address != cpu_instruction_master_address_last_time))
        begin
          $write("%0d ns: cpu_instruction_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_instruction_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_read_last_time <= 0;
      else 
        cpu_instruction_master_read_last_time <= cpu_instruction_master_read;
    end


  //cpu_instruction_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_instruction_master_read != cpu_instruction_master_read_last_time))
        begin
          $write("%0d ns: cpu_instruction_master_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_tightly_coupled_data_master_0_arbitrator (
                                                      // inputs:
                                                       clk,
                                                       cpu_tightly_coupled_data_master_0_address,
                                                       cpu_tightly_coupled_data_master_0_byteenable,
                                                       cpu_tightly_coupled_data_master_0_clken,
                                                       cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2,
                                                       cpu_tightly_coupled_data_master_0_qualified_request_tlb_miss_ram_1k_s2,
                                                       cpu_tightly_coupled_data_master_0_read,
                                                       cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2,
                                                       cpu_tightly_coupled_data_master_0_requests_tlb_miss_ram_1k_s2,
                                                       cpu_tightly_coupled_data_master_0_write,
                                                       cpu_tightly_coupled_data_master_0_writedata,
                                                       d1_tlb_miss_ram_1k_s2_end_xfer,
                                                       reset_n,
                                                       tlb_miss_ram_1k_s2_readdata_from_sa,

                                                      // outputs:
                                                       cpu_tightly_coupled_data_master_0_address_to_slave,
                                                       cpu_tightly_coupled_data_master_0_latency_counter,
                                                       cpu_tightly_coupled_data_master_0_readdata,
                                                       cpu_tightly_coupled_data_master_0_readdatavalid,
                                                       cpu_tightly_coupled_data_master_0_waitrequest
                                                    )
;

  output  [ 26: 0] cpu_tightly_coupled_data_master_0_address_to_slave;
  output           cpu_tightly_coupled_data_master_0_latency_counter;
  output  [ 31: 0] cpu_tightly_coupled_data_master_0_readdata;
  output           cpu_tightly_coupled_data_master_0_readdatavalid;
  output           cpu_tightly_coupled_data_master_0_waitrequest;
  input            clk;
  input   [ 26: 0] cpu_tightly_coupled_data_master_0_address;
  input   [  3: 0] cpu_tightly_coupled_data_master_0_byteenable;
  input            cpu_tightly_coupled_data_master_0_clken;
  input            cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2;
  input            cpu_tightly_coupled_data_master_0_qualified_request_tlb_miss_ram_1k_s2;
  input            cpu_tightly_coupled_data_master_0_read;
  input            cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2;
  input            cpu_tightly_coupled_data_master_0_requests_tlb_miss_ram_1k_s2;
  input            cpu_tightly_coupled_data_master_0_write;
  input   [ 31: 0] cpu_tightly_coupled_data_master_0_writedata;
  input            d1_tlb_miss_ram_1k_s2_end_xfer;
  input            reset_n;
  input   [ 31: 0] tlb_miss_ram_1k_s2_readdata_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 26: 0] cpu_tightly_coupled_data_master_0_address_last_time;
  wire    [ 26: 0] cpu_tightly_coupled_data_master_0_address_to_slave;
  reg     [  3: 0] cpu_tightly_coupled_data_master_0_byteenable_last_time;
  wire             cpu_tightly_coupled_data_master_0_latency_counter;
  reg              cpu_tightly_coupled_data_master_0_read_last_time;
  wire    [ 31: 0] cpu_tightly_coupled_data_master_0_readdata;
  wire             cpu_tightly_coupled_data_master_0_readdatavalid;
  wire             cpu_tightly_coupled_data_master_0_run;
  wire             cpu_tightly_coupled_data_master_0_waitrequest;
  reg              cpu_tightly_coupled_data_master_0_write_last_time;
  reg     [ 31: 0] cpu_tightly_coupled_data_master_0_writedata_last_time;
  wire             pre_flush_cpu_tightly_coupled_data_master_0_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & ((~cpu_tightly_coupled_data_master_0_qualified_request_tlb_miss_ram_1k_s2 | ~(cpu_tightly_coupled_data_master_0_read | cpu_tightly_coupled_data_master_0_write) | (1 & (cpu_tightly_coupled_data_master_0_read | cpu_tightly_coupled_data_master_0_write)))) & ((~cpu_tightly_coupled_data_master_0_qualified_request_tlb_miss_ram_1k_s2 | ~(cpu_tightly_coupled_data_master_0_read | cpu_tightly_coupled_data_master_0_write) | (1 & (cpu_tightly_coupled_data_master_0_read | cpu_tightly_coupled_data_master_0_write))));

  //cascaded wait assignment, which is an e_assign
  assign cpu_tightly_coupled_data_master_0_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_tightly_coupled_data_master_0_address_to_slave = {17'b11111111111111101,
    cpu_tightly_coupled_data_master_0_address[9 : 0]};

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_tightly_coupled_data_master_0_readdatavalid = cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_tightly_coupled_data_master_0_readdatavalid = 0 |
    pre_flush_cpu_tightly_coupled_data_master_0_readdatavalid;

  //cpu/tightly_coupled_data_master_0 readdata mux, which is an e_mux
  assign cpu_tightly_coupled_data_master_0_readdata = tlb_miss_ram_1k_s2_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign cpu_tightly_coupled_data_master_0_waitrequest = ~cpu_tightly_coupled_data_master_0_run;

  //latent max counter, which is an e_assign
  assign cpu_tightly_coupled_data_master_0_latency_counter = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_tightly_coupled_data_master_0_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_tightly_coupled_data_master_0_address_last_time <= 0;
      else 
        cpu_tightly_coupled_data_master_0_address_last_time <= cpu_tightly_coupled_data_master_0_address;
    end


  //cpu/tightly_coupled_data_master_0 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_tightly_coupled_data_master_0_waitrequest & (cpu_tightly_coupled_data_master_0_read | cpu_tightly_coupled_data_master_0_write);
    end


  //cpu_tightly_coupled_data_master_0_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_tightly_coupled_data_master_0_address != cpu_tightly_coupled_data_master_0_address_last_time))
        begin
          $write("%0d ns: cpu_tightly_coupled_data_master_0_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_tightly_coupled_data_master_0_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_tightly_coupled_data_master_0_byteenable_last_time <= 0;
      else 
        cpu_tightly_coupled_data_master_0_byteenable_last_time <= cpu_tightly_coupled_data_master_0_byteenable;
    end


  //cpu_tightly_coupled_data_master_0_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_tightly_coupled_data_master_0_byteenable != cpu_tightly_coupled_data_master_0_byteenable_last_time))
        begin
          $write("%0d ns: cpu_tightly_coupled_data_master_0_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_tightly_coupled_data_master_0_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_tightly_coupled_data_master_0_read_last_time <= 0;
      else 
        cpu_tightly_coupled_data_master_0_read_last_time <= cpu_tightly_coupled_data_master_0_read;
    end


  //cpu_tightly_coupled_data_master_0_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_tightly_coupled_data_master_0_read != cpu_tightly_coupled_data_master_0_read_last_time))
        begin
          $write("%0d ns: cpu_tightly_coupled_data_master_0_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_tightly_coupled_data_master_0_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_tightly_coupled_data_master_0_write_last_time <= 0;
      else 
        cpu_tightly_coupled_data_master_0_write_last_time <= cpu_tightly_coupled_data_master_0_write;
    end


  //cpu_tightly_coupled_data_master_0_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_tightly_coupled_data_master_0_write != cpu_tightly_coupled_data_master_0_write_last_time))
        begin
          $write("%0d ns: cpu_tightly_coupled_data_master_0_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_tightly_coupled_data_master_0_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_tightly_coupled_data_master_0_writedata_last_time <= 0;
      else 
        cpu_tightly_coupled_data_master_0_writedata_last_time <= cpu_tightly_coupled_data_master_0_writedata;
    end


  //cpu_tightly_coupled_data_master_0_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_tightly_coupled_data_master_0_writedata != cpu_tightly_coupled_data_master_0_writedata_last_time) & cpu_tightly_coupled_data_master_0_write)
        begin
          $write("%0d ns: cpu_tightly_coupled_data_master_0_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_tightly_coupled_instruction_master_0_arbitrator (
                                                             // inputs:
                                                              clk,
                                                              cpu_tightly_coupled_instruction_master_0_address,
                                                              cpu_tightly_coupled_instruction_master_0_clken,
                                                              cpu_tightly_coupled_instruction_master_0_granted_tlb_miss_ram_1k_s1,
                                                              cpu_tightly_coupled_instruction_master_0_qualified_request_tlb_miss_ram_1k_s1,
                                                              cpu_tightly_coupled_instruction_master_0_read,
                                                              cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1,
                                                              cpu_tightly_coupled_instruction_master_0_requests_tlb_miss_ram_1k_s1,
                                                              d1_tlb_miss_ram_1k_s1_end_xfer,
                                                              reset_n,
                                                              tlb_miss_ram_1k_s1_readdata_from_sa,

                                                             // outputs:
                                                              cpu_tightly_coupled_instruction_master_0_address_to_slave,
                                                              cpu_tightly_coupled_instruction_master_0_latency_counter,
                                                              cpu_tightly_coupled_instruction_master_0_readdata,
                                                              cpu_tightly_coupled_instruction_master_0_readdatavalid,
                                                              cpu_tightly_coupled_instruction_master_0_waitrequest
                                                           )
;

  output  [ 26: 0] cpu_tightly_coupled_instruction_master_0_address_to_slave;
  output           cpu_tightly_coupled_instruction_master_0_latency_counter;
  output  [ 31: 0] cpu_tightly_coupled_instruction_master_0_readdata;
  output           cpu_tightly_coupled_instruction_master_0_readdatavalid;
  output           cpu_tightly_coupled_instruction_master_0_waitrequest;
  input            clk;
  input   [ 26: 0] cpu_tightly_coupled_instruction_master_0_address;
  input            cpu_tightly_coupled_instruction_master_0_clken;
  input            cpu_tightly_coupled_instruction_master_0_granted_tlb_miss_ram_1k_s1;
  input            cpu_tightly_coupled_instruction_master_0_qualified_request_tlb_miss_ram_1k_s1;
  input            cpu_tightly_coupled_instruction_master_0_read;
  input            cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1;
  input            cpu_tightly_coupled_instruction_master_0_requests_tlb_miss_ram_1k_s1;
  input            d1_tlb_miss_ram_1k_s1_end_xfer;
  input            reset_n;
  input   [ 31: 0] tlb_miss_ram_1k_s1_readdata_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 26: 0] cpu_tightly_coupled_instruction_master_0_address_last_time;
  wire    [ 26: 0] cpu_tightly_coupled_instruction_master_0_address_to_slave;
  wire             cpu_tightly_coupled_instruction_master_0_latency_counter;
  reg              cpu_tightly_coupled_instruction_master_0_read_last_time;
  wire    [ 31: 0] cpu_tightly_coupled_instruction_master_0_readdata;
  wire             cpu_tightly_coupled_instruction_master_0_readdatavalid;
  wire             cpu_tightly_coupled_instruction_master_0_run;
  wire             cpu_tightly_coupled_instruction_master_0_waitrequest;
  wire             pre_flush_cpu_tightly_coupled_instruction_master_0_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & ((~cpu_tightly_coupled_instruction_master_0_qualified_request_tlb_miss_ram_1k_s1 | ~(cpu_tightly_coupled_instruction_master_0_read) | (1 & (cpu_tightly_coupled_instruction_master_0_read))));

  //cascaded wait assignment, which is an e_assign
  assign cpu_tightly_coupled_instruction_master_0_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_tightly_coupled_instruction_master_0_address_to_slave = {17'b11111111111111101,
    cpu_tightly_coupled_instruction_master_0_address[9 : 0]};

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_tightly_coupled_instruction_master_0_readdatavalid = cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_tightly_coupled_instruction_master_0_readdatavalid = 0 |
    pre_flush_cpu_tightly_coupled_instruction_master_0_readdatavalid;

  //cpu/tightly_coupled_instruction_master_0 readdata mux, which is an e_mux
  assign cpu_tightly_coupled_instruction_master_0_readdata = tlb_miss_ram_1k_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign cpu_tightly_coupled_instruction_master_0_waitrequest = ~cpu_tightly_coupled_instruction_master_0_run;

  //latent max counter, which is an e_assign
  assign cpu_tightly_coupled_instruction_master_0_latency_counter = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_tightly_coupled_instruction_master_0_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_tightly_coupled_instruction_master_0_address_last_time <= 0;
      else 
        cpu_tightly_coupled_instruction_master_0_address_last_time <= cpu_tightly_coupled_instruction_master_0_address;
    end


  //cpu/tightly_coupled_instruction_master_0 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_tightly_coupled_instruction_master_0_waitrequest & (cpu_tightly_coupled_instruction_master_0_read);
    end


  //cpu_tightly_coupled_instruction_master_0_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_tightly_coupled_instruction_master_0_address != cpu_tightly_coupled_instruction_master_0_address_last_time))
        begin
          $write("%0d ns: cpu_tightly_coupled_instruction_master_0_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_tightly_coupled_instruction_master_0_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_tightly_coupled_instruction_master_0_read_last_time <= 0;
      else 
        cpu_tightly_coupled_instruction_master_0_read_last_time <= cpu_tightly_coupled_instruction_master_0_read;
    end


  //cpu_tightly_coupled_instruction_master_0_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_tightly_coupled_instruction_master_0_read != cpu_tightly_coupled_instruction_master_0_read_last_time))
        begin
          $write("%0d ns: cpu_tightly_coupled_instruction_master_0_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_pb_cpu_to_ddr3_top_m1_to_ddr3_top_s1_module (
                                                                  // inputs:
                                                                   clear_fifo,
                                                                   clk,
                                                                   data_in,
                                                                   read,
                                                                   reset_n,
                                                                   sync_reset,
                                                                   write,

                                                                  // outputs:
                                                                   data_out,
                                                                   empty,
                                                                   fifo_contains_ones_n,
                                                                   full
                                                                )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  wire             full_32;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_31;
  assign empty = !full_0;
  assign full_32 = 0;
  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    0;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_pb_dma_to_ddr3_top_m1_to_ddr3_top_s1_module (
                                                                  // inputs:
                                                                   clear_fifo,
                                                                   clk,
                                                                   data_in,
                                                                   read,
                                                                   reset_n,
                                                                   sync_reset,
                                                                   write,

                                                                  // outputs:
                                                                   data_out,
                                                                   empty,
                                                                   fifo_contains_ones_n,
                                                                   full
                                                                )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  wire             full_32;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_31;
  assign empty = !full_0;
  assign full_32 = 0;
  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    0;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ddr3_top_s1_arbitrator (
                                // inputs:
                                 clk,
                                 ddr3_top_s1_readdata,
                                 ddr3_top_s1_readdatavalid,
                                 ddr3_top_s1_resetrequest_n,
                                 ddr3_top_s1_waitrequest_n,
                                 pb_cpu_to_ddr3_top_m1_address_to_slave,
                                 pb_cpu_to_ddr3_top_m1_burstcount,
                                 pb_cpu_to_ddr3_top_m1_byteenable,
                                 pb_cpu_to_ddr3_top_m1_chipselect,
                                 pb_cpu_to_ddr3_top_m1_latency_counter,
                                 pb_cpu_to_ddr3_top_m1_read,
                                 pb_cpu_to_ddr3_top_m1_write,
                                 pb_cpu_to_ddr3_top_m1_writedata,
                                 pb_dma_to_ddr3_top_m1_address_to_slave,
                                 pb_dma_to_ddr3_top_m1_burstcount,
                                 pb_dma_to_ddr3_top_m1_byteenable,
                                 pb_dma_to_ddr3_top_m1_chipselect,
                                 pb_dma_to_ddr3_top_m1_latency_counter,
                                 pb_dma_to_ddr3_top_m1_read,
                                 pb_dma_to_ddr3_top_m1_write,
                                 pb_dma_to_ddr3_top_m1_writedata,
                                 reset_n,

                                // outputs:
                                 d1_ddr3_top_s1_end_xfer,
                                 ddr3_top_s1_address,
                                 ddr3_top_s1_beginbursttransfer,
                                 ddr3_top_s1_burstcount,
                                 ddr3_top_s1_byteenable,
                                 ddr3_top_s1_read,
                                 ddr3_top_s1_readdata_from_sa,
                                 ddr3_top_s1_resetrequest_n_from_sa,
                                 ddr3_top_s1_waitrequest_n_from_sa,
                                 ddr3_top_s1_write,
                                 ddr3_top_s1_writedata,
                                 pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1,
                                 pb_cpu_to_ddr3_top_m1_qualified_request_ddr3_top_s1,
                                 pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1,
                                 pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register,
                                 pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1,
                                 pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1,
                                 pb_dma_to_ddr3_top_m1_qualified_request_ddr3_top_s1,
                                 pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1,
                                 pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register,
                                 pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1
                              )
;

  output           d1_ddr3_top_s1_end_xfer;
  output  [ 23: 0] ddr3_top_s1_address;
  output           ddr3_top_s1_beginbursttransfer;
  output  [  2: 0] ddr3_top_s1_burstcount;
  output  [  7: 0] ddr3_top_s1_byteenable;
  output           ddr3_top_s1_read;
  output  [ 63: 0] ddr3_top_s1_readdata_from_sa;
  output           ddr3_top_s1_resetrequest_n_from_sa;
  output           ddr3_top_s1_waitrequest_n_from_sa;
  output           ddr3_top_s1_write;
  output  [ 63: 0] ddr3_top_s1_writedata;
  output           pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1;
  output           pb_cpu_to_ddr3_top_m1_qualified_request_ddr3_top_s1;
  output           pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1;
  output           pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register;
  output           pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1;
  output           pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1;
  output           pb_dma_to_ddr3_top_m1_qualified_request_ddr3_top_s1;
  output           pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1;
  output           pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register;
  output           pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1;
  input            clk;
  input   [ 63: 0] ddr3_top_s1_readdata;
  input            ddr3_top_s1_readdatavalid;
  input            ddr3_top_s1_resetrequest_n;
  input            ddr3_top_s1_waitrequest_n;
  input   [ 26: 0] pb_cpu_to_ddr3_top_m1_address_to_slave;
  input            pb_cpu_to_ddr3_top_m1_burstcount;
  input   [  3: 0] pb_cpu_to_ddr3_top_m1_byteenable;
  input            pb_cpu_to_ddr3_top_m1_chipselect;
  input            pb_cpu_to_ddr3_top_m1_latency_counter;
  input            pb_cpu_to_ddr3_top_m1_read;
  input            pb_cpu_to_ddr3_top_m1_write;
  input   [ 31: 0] pb_cpu_to_ddr3_top_m1_writedata;
  input   [ 26: 0] pb_dma_to_ddr3_top_m1_address_to_slave;
  input            pb_dma_to_ddr3_top_m1_burstcount;
  input   [  3: 0] pb_dma_to_ddr3_top_m1_byteenable;
  input            pb_dma_to_ddr3_top_m1_chipselect;
  input            pb_dma_to_ddr3_top_m1_latency_counter;
  input            pb_dma_to_ddr3_top_m1_read;
  input            pb_dma_to_ddr3_top_m1_write;
  input   [ 31: 0] pb_dma_to_ddr3_top_m1_writedata;
  input            reset_n;

  reg              d1_ddr3_top_s1_end_xfer;
  reg              d1_reasons_to_wait;
  wire    [ 23: 0] ddr3_top_s1_address;
  wire             ddr3_top_s1_allgrants;
  wire             ddr3_top_s1_allow_new_arb_cycle;
  wire             ddr3_top_s1_any_bursting_master_saved_grant;
  wire             ddr3_top_s1_any_continuerequest;
  reg     [  1: 0] ddr3_top_s1_arb_addend;
  wire             ddr3_top_s1_arb_counter_enable;
  reg     [  3: 0] ddr3_top_s1_arb_share_counter;
  wire    [  3: 0] ddr3_top_s1_arb_share_counter_next_value;
  wire    [  3: 0] ddr3_top_s1_arb_share_set_values;
  wire    [  1: 0] ddr3_top_s1_arb_winner;
  wire             ddr3_top_s1_arbitration_holdoff_internal;
  reg     [  1: 0] ddr3_top_s1_bbt_burstcounter;
  wire             ddr3_top_s1_beginbursttransfer;
  wire             ddr3_top_s1_beginbursttransfer_internal;
  wire             ddr3_top_s1_begins_xfer;
  wire    [  2: 0] ddr3_top_s1_burstcount;
  wire    [  7: 0] ddr3_top_s1_byteenable;
  wire    [  3: 0] ddr3_top_s1_chosen_master_double_vector;
  wire    [  1: 0] ddr3_top_s1_chosen_master_rot_left;
  wire             ddr3_top_s1_end_xfer;
  wire             ddr3_top_s1_firsttransfer;
  wire    [  1: 0] ddr3_top_s1_grant_vector;
  wire             ddr3_top_s1_in_a_read_cycle;
  wire             ddr3_top_s1_in_a_write_cycle;
  wire    [  1: 0] ddr3_top_s1_master_qreq_vector;
  wire             ddr3_top_s1_move_on_to_next_transaction;
  wire    [  1: 0] ddr3_top_s1_next_bbt_burstcount;
  wire             ddr3_top_s1_non_bursting_master_requests;
  wire             ddr3_top_s1_read;
  wire    [ 63: 0] ddr3_top_s1_readdata_from_sa;
  wire             ddr3_top_s1_readdatavalid_from_sa;
  reg              ddr3_top_s1_reg_firsttransfer;
  wire             ddr3_top_s1_resetrequest_n_from_sa;
  reg     [  1: 0] ddr3_top_s1_saved_chosen_master_vector;
  reg              ddr3_top_s1_slavearbiterlockenable;
  wire             ddr3_top_s1_slavearbiterlockenable2;
  wire             ddr3_top_s1_unreg_firsttransfer;
  wire             ddr3_top_s1_waitrequest_n_from_sa;
  wire             ddr3_top_s1_waits_for_read;
  wire             ddr3_top_s1_waits_for_write;
  wire             ddr3_top_s1_write;
  wire    [ 63: 0] ddr3_top_s1_writedata;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_ddr3_top_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_pb_cpu_to_ddr3_top_m1_granted_slave_ddr3_top_s1;
  reg              last_cycle_pb_dma_to_ddr3_top_m1_granted_slave_ddr3_top_s1;
  wire             pb_cpu_to_ddr3_top_m1_arbiterlock;
  wire             pb_cpu_to_ddr3_top_m1_arbiterlock2;
  wire    [  7: 0] pb_cpu_to_ddr3_top_m1_byteenable_ddr3_top_s1;
  wire             pb_cpu_to_ddr3_top_m1_continuerequest;
  wire             pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1;
  wire             pb_cpu_to_ddr3_top_m1_qualified_request_ddr3_top_s1;
  wire             pb_cpu_to_ddr3_top_m1_rdv_fifo_empty_ddr3_top_s1;
  wire             pb_cpu_to_ddr3_top_m1_rdv_fifo_output_from_ddr3_top_s1;
  wire             pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1;
  wire             pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register;
  wire             pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1;
  wire             pb_cpu_to_ddr3_top_m1_saved_grant_ddr3_top_s1;
  wire    [ 63: 0] pb_cpu_to_ddr3_top_m1_writedata_replicated;
  wire             pb_dma_to_ddr3_top_m1_arbiterlock;
  wire             pb_dma_to_ddr3_top_m1_arbiterlock2;
  wire    [  7: 0] pb_dma_to_ddr3_top_m1_byteenable_ddr3_top_s1;
  wire             pb_dma_to_ddr3_top_m1_continuerequest;
  wire             pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1;
  wire             pb_dma_to_ddr3_top_m1_qualified_request_ddr3_top_s1;
  wire             pb_dma_to_ddr3_top_m1_rdv_fifo_empty_ddr3_top_s1;
  wire             pb_dma_to_ddr3_top_m1_rdv_fifo_output_from_ddr3_top_s1;
  wire             pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1;
  wire             pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register;
  wire             pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1;
  wire             pb_dma_to_ddr3_top_m1_saved_grant_ddr3_top_s1;
  wire    [ 63: 0] pb_dma_to_ddr3_top_m1_writedata_replicated;
  wire    [ 26: 0] shifted_address_to_ddr3_top_s1_from_pb_cpu_to_ddr3_top_m1;
  wire    [ 26: 0] shifted_address_to_ddr3_top_s1_from_pb_dma_to_ddr3_top_m1;
  wire             wait_for_ddr3_top_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~ddr3_top_s1_end_xfer;
    end


  assign ddr3_top_s1_begins_xfer = ~d1_reasons_to_wait & ((pb_cpu_to_ddr3_top_m1_qualified_request_ddr3_top_s1 | pb_dma_to_ddr3_top_m1_qualified_request_ddr3_top_s1));
  //assign ddr3_top_s1_readdata_from_sa = ddr3_top_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr3_top_s1_readdata_from_sa = ddr3_top_s1_readdata;

  assign pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1 = (1) & pb_cpu_to_ddr3_top_m1_chipselect;
  //assign ddr3_top_s1_waitrequest_n_from_sa = ddr3_top_s1_waitrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr3_top_s1_waitrequest_n_from_sa = ddr3_top_s1_waitrequest_n;

  //assign ddr3_top_s1_readdatavalid_from_sa = ddr3_top_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr3_top_s1_readdatavalid_from_sa = ddr3_top_s1_readdatavalid;

  //ddr3_top_s1_arb_share_counter set values, which is an e_mux
  assign ddr3_top_s1_arb_share_set_values = (pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1)? 8 :
    (pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1)? 8 :
    (pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1)? 8 :
    (pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1)? 8 :
    1;

  //ddr3_top_s1_non_bursting_master_requests mux, which is an e_mux
  assign ddr3_top_s1_non_bursting_master_requests = pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1 |
    pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1 |
    pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1 |
    pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1;

  //ddr3_top_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign ddr3_top_s1_any_bursting_master_saved_grant = 0;

  //ddr3_top_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign ddr3_top_s1_arb_share_counter_next_value = ddr3_top_s1_firsttransfer ? (ddr3_top_s1_arb_share_set_values - 1) : |ddr3_top_s1_arb_share_counter ? (ddr3_top_s1_arb_share_counter - 1) : 0;

  //ddr3_top_s1_allgrants all slave grants, which is an e_mux
  assign ddr3_top_s1_allgrants = (|ddr3_top_s1_grant_vector) |
    (|ddr3_top_s1_grant_vector) |
    (|ddr3_top_s1_grant_vector) |
    (|ddr3_top_s1_grant_vector);

  //ddr3_top_s1_end_xfer assignment, which is an e_assign
  assign ddr3_top_s1_end_xfer = ~(ddr3_top_s1_waits_for_read | ddr3_top_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_ddr3_top_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_ddr3_top_s1 = ddr3_top_s1_end_xfer & (~ddr3_top_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //ddr3_top_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign ddr3_top_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_ddr3_top_s1 & ddr3_top_s1_allgrants) | (end_xfer_arb_share_counter_term_ddr3_top_s1 & ~ddr3_top_s1_non_bursting_master_requests);

  //ddr3_top_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr3_top_s1_arb_share_counter <= 0;
      else if (ddr3_top_s1_arb_counter_enable)
          ddr3_top_s1_arb_share_counter <= ddr3_top_s1_arb_share_counter_next_value;
    end


  //ddr3_top_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr3_top_s1_slavearbiterlockenable <= 0;
      else if ((|ddr3_top_s1_master_qreq_vector & end_xfer_arb_share_counter_term_ddr3_top_s1) | (end_xfer_arb_share_counter_term_ddr3_top_s1 & ~ddr3_top_s1_non_bursting_master_requests))
          ddr3_top_s1_slavearbiterlockenable <= |ddr3_top_s1_arb_share_counter_next_value;
    end


  //pb_cpu_to_ddr3_top/m1 ddr3_top/s1 arbiterlock, which is an e_assign
  assign pb_cpu_to_ddr3_top_m1_arbiterlock = ddr3_top_s1_slavearbiterlockenable & pb_cpu_to_ddr3_top_m1_continuerequest;

  //ddr3_top_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign ddr3_top_s1_slavearbiterlockenable2 = |ddr3_top_s1_arb_share_counter_next_value;

  //pb_cpu_to_ddr3_top/m1 ddr3_top/s1 arbiterlock2, which is an e_assign
  assign pb_cpu_to_ddr3_top_m1_arbiterlock2 = ddr3_top_s1_slavearbiterlockenable2 & pb_cpu_to_ddr3_top_m1_continuerequest;

  //pb_dma_to_ddr3_top/m1 ddr3_top/s1 arbiterlock, which is an e_assign
  assign pb_dma_to_ddr3_top_m1_arbiterlock = ddr3_top_s1_slavearbiterlockenable & pb_dma_to_ddr3_top_m1_continuerequest;

  //pb_dma_to_ddr3_top/m1 ddr3_top/s1 arbiterlock2, which is an e_assign
  assign pb_dma_to_ddr3_top_m1_arbiterlock2 = ddr3_top_s1_slavearbiterlockenable2 & pb_dma_to_ddr3_top_m1_continuerequest;

  //pb_dma_to_ddr3_top/m1 granted ddr3_top/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_pb_dma_to_ddr3_top_m1_granted_slave_ddr3_top_s1 <= 0;
      else 
        last_cycle_pb_dma_to_ddr3_top_m1_granted_slave_ddr3_top_s1 <= pb_dma_to_ddr3_top_m1_saved_grant_ddr3_top_s1 ? 1 : (ddr3_top_s1_arbitration_holdoff_internal | ~pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1) ? 0 : last_cycle_pb_dma_to_ddr3_top_m1_granted_slave_ddr3_top_s1;
    end


  //pb_dma_to_ddr3_top_m1_continuerequest continued request, which is an e_mux
  assign pb_dma_to_ddr3_top_m1_continuerequest = last_cycle_pb_dma_to_ddr3_top_m1_granted_slave_ddr3_top_s1 & pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1;

  //ddr3_top_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign ddr3_top_s1_any_continuerequest = pb_dma_to_ddr3_top_m1_continuerequest |
    pb_cpu_to_ddr3_top_m1_continuerequest;

  assign pb_cpu_to_ddr3_top_m1_qualified_request_ddr3_top_s1 = pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1 & ~(((pb_cpu_to_ddr3_top_m1_read & pb_cpu_to_ddr3_top_m1_chipselect) & ((pb_cpu_to_ddr3_top_m1_latency_counter != 0) | (1 < pb_cpu_to_ddr3_top_m1_latency_counter))) | pb_dma_to_ddr3_top_m1_arbiterlock);
  //unique name for ddr3_top_s1_move_on_to_next_transaction, which is an e_assign
  assign ddr3_top_s1_move_on_to_next_transaction = ddr3_top_s1_readdatavalid_from_sa;

  //rdv_fifo_for_pb_cpu_to_ddr3_top_m1_to_ddr3_top_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_pb_cpu_to_ddr3_top_m1_to_ddr3_top_s1_module rdv_fifo_for_pb_cpu_to_ddr3_top_m1_to_ddr3_top_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1),
      .data_out             (pb_cpu_to_ddr3_top_m1_rdv_fifo_output_from_ddr3_top_s1),
      .empty                (),
      .fifo_contains_ones_n (pb_cpu_to_ddr3_top_m1_rdv_fifo_empty_ddr3_top_s1),
      .full                 (),
      .read                 (ddr3_top_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~ddr3_top_s1_waits_for_read)
    );

  assign pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register = ~pb_cpu_to_ddr3_top_m1_rdv_fifo_empty_ddr3_top_s1;
  //local readdatavalid pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1, which is an e_mux
  assign pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1 = (ddr3_top_s1_readdatavalid_from_sa & pb_cpu_to_ddr3_top_m1_rdv_fifo_output_from_ddr3_top_s1) & ~ pb_cpu_to_ddr3_top_m1_rdv_fifo_empty_ddr3_top_s1;

  //replicate narrow data for wide slave
  assign pb_cpu_to_ddr3_top_m1_writedata_replicated = {pb_cpu_to_ddr3_top_m1_writedata,
    pb_cpu_to_ddr3_top_m1_writedata};

  //ddr3_top_s1_writedata mux, which is an e_mux
  assign ddr3_top_s1_writedata = (pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1)? pb_cpu_to_ddr3_top_m1_writedata_replicated :
    pb_dma_to_ddr3_top_m1_writedata_replicated;

  assign pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1 = (1) & pb_dma_to_ddr3_top_m1_chipselect;
  //pb_cpu_to_ddr3_top/m1 granted ddr3_top/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_pb_cpu_to_ddr3_top_m1_granted_slave_ddr3_top_s1 <= 0;
      else 
        last_cycle_pb_cpu_to_ddr3_top_m1_granted_slave_ddr3_top_s1 <= pb_cpu_to_ddr3_top_m1_saved_grant_ddr3_top_s1 ? 1 : (ddr3_top_s1_arbitration_holdoff_internal | ~pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1) ? 0 : last_cycle_pb_cpu_to_ddr3_top_m1_granted_slave_ddr3_top_s1;
    end


  //pb_cpu_to_ddr3_top_m1_continuerequest continued request, which is an e_mux
  assign pb_cpu_to_ddr3_top_m1_continuerequest = last_cycle_pb_cpu_to_ddr3_top_m1_granted_slave_ddr3_top_s1 & pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1;

  assign pb_dma_to_ddr3_top_m1_qualified_request_ddr3_top_s1 = pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1 & ~(((pb_dma_to_ddr3_top_m1_read & pb_dma_to_ddr3_top_m1_chipselect) & ((pb_dma_to_ddr3_top_m1_latency_counter != 0) | (1 < pb_dma_to_ddr3_top_m1_latency_counter))) | pb_cpu_to_ddr3_top_m1_arbiterlock);
  //rdv_fifo_for_pb_dma_to_ddr3_top_m1_to_ddr3_top_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_pb_dma_to_ddr3_top_m1_to_ddr3_top_s1_module rdv_fifo_for_pb_dma_to_ddr3_top_m1_to_ddr3_top_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1),
      .data_out             (pb_dma_to_ddr3_top_m1_rdv_fifo_output_from_ddr3_top_s1),
      .empty                (),
      .fifo_contains_ones_n (pb_dma_to_ddr3_top_m1_rdv_fifo_empty_ddr3_top_s1),
      .full                 (),
      .read                 (ddr3_top_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~ddr3_top_s1_waits_for_read)
    );

  assign pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register = ~pb_dma_to_ddr3_top_m1_rdv_fifo_empty_ddr3_top_s1;
  //local readdatavalid pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1, which is an e_mux
  assign pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1 = (ddr3_top_s1_readdatavalid_from_sa & pb_dma_to_ddr3_top_m1_rdv_fifo_output_from_ddr3_top_s1) & ~ pb_dma_to_ddr3_top_m1_rdv_fifo_empty_ddr3_top_s1;

  //replicate narrow data for wide slave
  assign pb_dma_to_ddr3_top_m1_writedata_replicated = {pb_dma_to_ddr3_top_m1_writedata,
    pb_dma_to_ddr3_top_m1_writedata};

  //allow new arb cycle for ddr3_top/s1, which is an e_assign
  assign ddr3_top_s1_allow_new_arb_cycle = ~pb_cpu_to_ddr3_top_m1_arbiterlock & ~pb_dma_to_ddr3_top_m1_arbiterlock;

  //pb_dma_to_ddr3_top/m1 assignment into master qualified-requests vector for ddr3_top/s1, which is an e_assign
  assign ddr3_top_s1_master_qreq_vector[0] = pb_dma_to_ddr3_top_m1_qualified_request_ddr3_top_s1;

  //pb_dma_to_ddr3_top/m1 grant ddr3_top/s1, which is an e_assign
  assign pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1 = ddr3_top_s1_grant_vector[0];

  //pb_dma_to_ddr3_top/m1 saved-grant ddr3_top/s1, which is an e_assign
  assign pb_dma_to_ddr3_top_m1_saved_grant_ddr3_top_s1 = ddr3_top_s1_arb_winner[0] && pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1;

  //pb_cpu_to_ddr3_top/m1 assignment into master qualified-requests vector for ddr3_top/s1, which is an e_assign
  assign ddr3_top_s1_master_qreq_vector[1] = pb_cpu_to_ddr3_top_m1_qualified_request_ddr3_top_s1;

  //pb_cpu_to_ddr3_top/m1 grant ddr3_top/s1, which is an e_assign
  assign pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1 = ddr3_top_s1_grant_vector[1];

  //pb_cpu_to_ddr3_top/m1 saved-grant ddr3_top/s1, which is an e_assign
  assign pb_cpu_to_ddr3_top_m1_saved_grant_ddr3_top_s1 = ddr3_top_s1_arb_winner[1] && pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1;

  //ddr3_top/s1 chosen-master double-vector, which is an e_assign
  assign ddr3_top_s1_chosen_master_double_vector = {ddr3_top_s1_master_qreq_vector, ddr3_top_s1_master_qreq_vector} & ({~ddr3_top_s1_master_qreq_vector, ~ddr3_top_s1_master_qreq_vector} + ddr3_top_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign ddr3_top_s1_arb_winner = (ddr3_top_s1_allow_new_arb_cycle & | ddr3_top_s1_grant_vector) ? ddr3_top_s1_grant_vector : ddr3_top_s1_saved_chosen_master_vector;

  //saved ddr3_top_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr3_top_s1_saved_chosen_master_vector <= 0;
      else if (ddr3_top_s1_allow_new_arb_cycle)
          ddr3_top_s1_saved_chosen_master_vector <= |ddr3_top_s1_grant_vector ? ddr3_top_s1_grant_vector : ddr3_top_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign ddr3_top_s1_grant_vector = {(ddr3_top_s1_chosen_master_double_vector[1] | ddr3_top_s1_chosen_master_double_vector[3]),
    (ddr3_top_s1_chosen_master_double_vector[0] | ddr3_top_s1_chosen_master_double_vector[2])};

  //ddr3_top/s1 chosen master rotated left, which is an e_assign
  assign ddr3_top_s1_chosen_master_rot_left = (ddr3_top_s1_arb_winner << 1) ? (ddr3_top_s1_arb_winner << 1) : 1;

  //ddr3_top/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr3_top_s1_arb_addend <= 1;
      else if (|ddr3_top_s1_grant_vector)
          ddr3_top_s1_arb_addend <= ddr3_top_s1_end_xfer? ddr3_top_s1_chosen_master_rot_left : ddr3_top_s1_grant_vector;
    end


  //assign ddr3_top_s1_resetrequest_n_from_sa = ddr3_top_s1_resetrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr3_top_s1_resetrequest_n_from_sa = ddr3_top_s1_resetrequest_n;

  //ddr3_top_s1_firsttransfer first transaction, which is an e_assign
  assign ddr3_top_s1_firsttransfer = ddr3_top_s1_begins_xfer ? ddr3_top_s1_unreg_firsttransfer : ddr3_top_s1_reg_firsttransfer;

  //ddr3_top_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign ddr3_top_s1_unreg_firsttransfer = ~(ddr3_top_s1_slavearbiterlockenable & ddr3_top_s1_any_continuerequest);

  //ddr3_top_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr3_top_s1_reg_firsttransfer <= 1'b1;
      else if (ddr3_top_s1_begins_xfer)
          ddr3_top_s1_reg_firsttransfer <= ddr3_top_s1_unreg_firsttransfer;
    end


  //ddr3_top_s1_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign ddr3_top_s1_next_bbt_burstcount = ((((ddr3_top_s1_write) && (ddr3_top_s1_bbt_burstcounter == 0))))? (ddr3_top_s1_burstcount - 1) :
    ((((ddr3_top_s1_read) && (ddr3_top_s1_bbt_burstcounter == 0))))? 0 :
    (ddr3_top_s1_bbt_burstcounter - 1);

  //ddr3_top_s1_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr3_top_s1_bbt_burstcounter <= 0;
      else if (ddr3_top_s1_begins_xfer)
          ddr3_top_s1_bbt_burstcounter <= ddr3_top_s1_next_bbt_burstcount;
    end


  //ddr3_top_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign ddr3_top_s1_beginbursttransfer_internal = ddr3_top_s1_begins_xfer & (ddr3_top_s1_bbt_burstcounter == 0);

  //ddr3_top/s1 begin burst transfer to slave, which is an e_assign
  assign ddr3_top_s1_beginbursttransfer = ddr3_top_s1_beginbursttransfer_internal;

  //ddr3_top_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign ddr3_top_s1_arbitration_holdoff_internal = ddr3_top_s1_begins_xfer & ddr3_top_s1_firsttransfer;

  //ddr3_top_s1_read assignment, which is an e_mux
  assign ddr3_top_s1_read = (pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1 & (pb_cpu_to_ddr3_top_m1_read & pb_cpu_to_ddr3_top_m1_chipselect)) | (pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1 & (pb_dma_to_ddr3_top_m1_read & pb_dma_to_ddr3_top_m1_chipselect));

  //ddr3_top_s1_write assignment, which is an e_mux
  assign ddr3_top_s1_write = (pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1 & (pb_cpu_to_ddr3_top_m1_write & pb_cpu_to_ddr3_top_m1_chipselect)) | (pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1 & (pb_dma_to_ddr3_top_m1_write & pb_dma_to_ddr3_top_m1_chipselect));

  assign shifted_address_to_ddr3_top_s1_from_pb_cpu_to_ddr3_top_m1 = pb_cpu_to_ddr3_top_m1_address_to_slave;
  //ddr3_top_s1_address mux, which is an e_mux
  assign ddr3_top_s1_address = (pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1)? (shifted_address_to_ddr3_top_s1_from_pb_cpu_to_ddr3_top_m1 >> 3) :
    (shifted_address_to_ddr3_top_s1_from_pb_dma_to_ddr3_top_m1 >> 3);

  assign shifted_address_to_ddr3_top_s1_from_pb_dma_to_ddr3_top_m1 = pb_dma_to_ddr3_top_m1_address_to_slave;
  //d1_ddr3_top_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_ddr3_top_s1_end_xfer <= 1;
      else 
        d1_ddr3_top_s1_end_xfer <= ddr3_top_s1_end_xfer;
    end


  //ddr3_top_s1_waits_for_read in a cycle, which is an e_mux
  assign ddr3_top_s1_waits_for_read = ddr3_top_s1_in_a_read_cycle & ~ddr3_top_s1_waitrequest_n_from_sa;

  //ddr3_top_s1_in_a_read_cycle assignment, which is an e_assign
  assign ddr3_top_s1_in_a_read_cycle = (pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1 & (pb_cpu_to_ddr3_top_m1_read & pb_cpu_to_ddr3_top_m1_chipselect)) | (pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1 & (pb_dma_to_ddr3_top_m1_read & pb_dma_to_ddr3_top_m1_chipselect));

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = ddr3_top_s1_in_a_read_cycle;

  //ddr3_top_s1_waits_for_write in a cycle, which is an e_mux
  assign ddr3_top_s1_waits_for_write = ddr3_top_s1_in_a_write_cycle & ~ddr3_top_s1_waitrequest_n_from_sa;

  //ddr3_top_s1_in_a_write_cycle assignment, which is an e_assign
  assign ddr3_top_s1_in_a_write_cycle = (pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1 & (pb_cpu_to_ddr3_top_m1_write & pb_cpu_to_ddr3_top_m1_chipselect)) | (pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1 & (pb_dma_to_ddr3_top_m1_write & pb_dma_to_ddr3_top_m1_chipselect));

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = ddr3_top_s1_in_a_write_cycle;

  assign wait_for_ddr3_top_s1_counter = 0;
  //ddr3_top_s1_byteenable byte enable port mux, which is an e_mux
  assign ddr3_top_s1_byteenable = (pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1)? pb_cpu_to_ddr3_top_m1_byteenable_ddr3_top_s1 :
    (pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1)? pb_dma_to_ddr3_top_m1_byteenable_ddr3_top_s1 :
    -1;

  //byte_enable_mux for pb_cpu_to_ddr3_top/m1 and ddr3_top/s1, which is an e_mux
  assign pb_cpu_to_ddr3_top_m1_byteenable_ddr3_top_s1 = (pb_cpu_to_ddr3_top_m1_address_to_slave[2] == 0)? pb_cpu_to_ddr3_top_m1_byteenable :
    {pb_cpu_to_ddr3_top_m1_byteenable, {4'b0}};

  //byte_enable_mux for pb_dma_to_ddr3_top/m1 and ddr3_top/s1, which is an e_mux
  assign pb_dma_to_ddr3_top_m1_byteenable_ddr3_top_s1 = (pb_dma_to_ddr3_top_m1_address_to_slave[2] == 0)? pb_dma_to_ddr3_top_m1_byteenable :
    {pb_dma_to_ddr3_top_m1_byteenable, {4'b0}};

  //burstcount mux, which is an e_mux
  assign ddr3_top_s1_burstcount = (pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1)? pb_cpu_to_ddr3_top_m1_burstcount :
    (pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1)? pb_dma_to_ddr3_top_m1_burstcount :
    1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //ddr3_top/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pb_cpu_to_ddr3_top/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1 && (pb_cpu_to_ddr3_top_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pb_cpu_to_ddr3_top/m1 drove 0 on its 'burstcount' port while accessing slave ddr3_top/s1", $time);
          $stop;
        end
    end


  //pb_dma_to_ddr3_top/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1 && (pb_dma_to_ddr3_top_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pb_dma_to_ddr3_top/m1 drove 0 on its 'burstcount' port while accessing slave ddr3_top/s1", $time);
          $stop;
        end
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1 + pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_ddr3_top_m1_saved_grant_ddr3_top_s1 + pb_dma_to_ddr3_top_m1_saved_grant_ddr3_top_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ghrd_4sgx230_sopc_reset_clkin_100_domain_synch_module (
                                                               // inputs:
                                                                clk,
                                                                data_in,
                                                                reset_n,

                                                               // outputs:
                                                                data_out
                                                             )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module descriptor_memory_s1_arbitrator (
                                         // inputs:
                                          clk,
                                          descriptor_memory_s1_readdata,
                                          pb_cpu_to_io_m1_address_to_slave,
                                          pb_cpu_to_io_m1_burstcount,
                                          pb_cpu_to_io_m1_byteenable,
                                          pb_cpu_to_io_m1_chipselect,
                                          pb_cpu_to_io_m1_latency_counter,
                                          pb_cpu_to_io_m1_read,
                                          pb_cpu_to_io_m1_write,
                                          pb_cpu_to_io_m1_writedata,
                                          pb_dma_to_descriptor_memory_m1_address_to_slave,
                                          pb_dma_to_descriptor_memory_m1_burstcount,
                                          pb_dma_to_descriptor_memory_m1_byteenable,
                                          pb_dma_to_descriptor_memory_m1_chipselect,
                                          pb_dma_to_descriptor_memory_m1_latency_counter,
                                          pb_dma_to_descriptor_memory_m1_read,
                                          pb_dma_to_descriptor_memory_m1_write,
                                          pb_dma_to_descriptor_memory_m1_writedata,
                                          reset_n,

                                         // outputs:
                                          d1_descriptor_memory_s1_end_xfer,
                                          descriptor_memory_s1_address,
                                          descriptor_memory_s1_byteenable,
                                          descriptor_memory_s1_chipselect,
                                          descriptor_memory_s1_clken,
                                          descriptor_memory_s1_readdata_from_sa,
                                          descriptor_memory_s1_reset,
                                          descriptor_memory_s1_write,
                                          descriptor_memory_s1_writedata,
                                          pb_cpu_to_io_m1_granted_descriptor_memory_s1,
                                          pb_cpu_to_io_m1_qualified_request_descriptor_memory_s1,
                                          pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1,
                                          pb_cpu_to_io_m1_requests_descriptor_memory_s1,
                                          pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1,
                                          pb_dma_to_descriptor_memory_m1_qualified_request_descriptor_memory_s1,
                                          pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1,
                                          pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1
                                       )
;

  output           d1_descriptor_memory_s1_end_xfer;
  output  [ 10: 0] descriptor_memory_s1_address;
  output  [  3: 0] descriptor_memory_s1_byteenable;
  output           descriptor_memory_s1_chipselect;
  output           descriptor_memory_s1_clken;
  output  [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  output           descriptor_memory_s1_reset;
  output           descriptor_memory_s1_write;
  output  [ 31: 0] descriptor_memory_s1_writedata;
  output           pb_cpu_to_io_m1_granted_descriptor_memory_s1;
  output           pb_cpu_to_io_m1_qualified_request_descriptor_memory_s1;
  output           pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1;
  output           pb_cpu_to_io_m1_requests_descriptor_memory_s1;
  output           pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1;
  output           pb_dma_to_descriptor_memory_m1_qualified_request_descriptor_memory_s1;
  output           pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1;
  output           pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1;
  input            clk;
  input   [ 31: 0] descriptor_memory_s1_readdata;
  input   [ 22: 0] pb_cpu_to_io_m1_address_to_slave;
  input            pb_cpu_to_io_m1_burstcount;
  input   [  3: 0] pb_cpu_to_io_m1_byteenable;
  input            pb_cpu_to_io_m1_chipselect;
  input            pb_cpu_to_io_m1_latency_counter;
  input            pb_cpu_to_io_m1_read;
  input            pb_cpu_to_io_m1_write;
  input   [ 31: 0] pb_cpu_to_io_m1_writedata;
  input   [ 13: 0] pb_dma_to_descriptor_memory_m1_address_to_slave;
  input            pb_dma_to_descriptor_memory_m1_burstcount;
  input   [  3: 0] pb_dma_to_descriptor_memory_m1_byteenable;
  input            pb_dma_to_descriptor_memory_m1_chipselect;
  input            pb_dma_to_descriptor_memory_m1_latency_counter;
  input            pb_dma_to_descriptor_memory_m1_read;
  input            pb_dma_to_descriptor_memory_m1_write;
  input   [ 31: 0] pb_dma_to_descriptor_memory_m1_writedata;
  input            reset_n;

  reg              d1_descriptor_memory_s1_end_xfer;
  reg              d1_reasons_to_wait;
  wire    [ 10: 0] descriptor_memory_s1_address;
  wire             descriptor_memory_s1_allgrants;
  wire             descriptor_memory_s1_allow_new_arb_cycle;
  wire             descriptor_memory_s1_any_bursting_master_saved_grant;
  wire             descriptor_memory_s1_any_continuerequest;
  reg     [  1: 0] descriptor_memory_s1_arb_addend;
  wire             descriptor_memory_s1_arb_counter_enable;
  reg     [  3: 0] descriptor_memory_s1_arb_share_counter;
  wire    [  3: 0] descriptor_memory_s1_arb_share_counter_next_value;
  wire    [  3: 0] descriptor_memory_s1_arb_share_set_values;
  wire    [  1: 0] descriptor_memory_s1_arb_winner;
  wire             descriptor_memory_s1_arbitration_holdoff_internal;
  wire             descriptor_memory_s1_beginbursttransfer_internal;
  wire             descriptor_memory_s1_begins_xfer;
  wire    [  3: 0] descriptor_memory_s1_byteenable;
  wire             descriptor_memory_s1_chipselect;
  wire    [  3: 0] descriptor_memory_s1_chosen_master_double_vector;
  wire    [  1: 0] descriptor_memory_s1_chosen_master_rot_left;
  wire             descriptor_memory_s1_clken;
  wire             descriptor_memory_s1_end_xfer;
  wire             descriptor_memory_s1_firsttransfer;
  wire    [  1: 0] descriptor_memory_s1_grant_vector;
  wire             descriptor_memory_s1_in_a_read_cycle;
  wire             descriptor_memory_s1_in_a_write_cycle;
  wire    [  1: 0] descriptor_memory_s1_master_qreq_vector;
  wire             descriptor_memory_s1_non_bursting_master_requests;
  wire    [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  reg              descriptor_memory_s1_reg_firsttransfer;
  wire             descriptor_memory_s1_reset;
  reg     [  1: 0] descriptor_memory_s1_saved_chosen_master_vector;
  reg              descriptor_memory_s1_slavearbiterlockenable;
  wire             descriptor_memory_s1_slavearbiterlockenable2;
  wire             descriptor_memory_s1_unreg_firsttransfer;
  wire             descriptor_memory_s1_waits_for_read;
  wire             descriptor_memory_s1_waits_for_write;
  wire             descriptor_memory_s1_write;
  wire    [ 31: 0] descriptor_memory_s1_writedata;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_descriptor_memory_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_pb_cpu_to_io_m1_granted_slave_descriptor_memory_s1;
  reg              last_cycle_pb_dma_to_descriptor_memory_m1_granted_slave_descriptor_memory_s1;
  wire             p1_pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1_shift_register;
  wire             p1_pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1_shift_register;
  wire             pb_cpu_to_io_m1_arbiterlock;
  wire             pb_cpu_to_io_m1_arbiterlock2;
  wire             pb_cpu_to_io_m1_continuerequest;
  wire             pb_cpu_to_io_m1_granted_descriptor_memory_s1;
  wire             pb_cpu_to_io_m1_qualified_request_descriptor_memory_s1;
  wire             pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1;
  reg              pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1_shift_register;
  wire             pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1_shift_register_in;
  wire             pb_cpu_to_io_m1_requests_descriptor_memory_s1;
  wire             pb_cpu_to_io_m1_saved_grant_descriptor_memory_s1;
  wire             pb_dma_to_descriptor_memory_m1_arbiterlock;
  wire             pb_dma_to_descriptor_memory_m1_arbiterlock2;
  wire             pb_dma_to_descriptor_memory_m1_continuerequest;
  wire             pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1;
  wire             pb_dma_to_descriptor_memory_m1_qualified_request_descriptor_memory_s1;
  wire             pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1;
  reg              pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1_shift_register;
  wire             pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1_shift_register_in;
  wire             pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1;
  wire             pb_dma_to_descriptor_memory_m1_saved_grant_descriptor_memory_s1;
  wire    [ 22: 0] shifted_address_to_descriptor_memory_s1_from_pb_cpu_to_io_m1;
  wire    [ 13: 0] shifted_address_to_descriptor_memory_s1_from_pb_dma_to_descriptor_memory_m1;
  wire             wait_for_descriptor_memory_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~descriptor_memory_s1_end_xfer;
    end


  assign descriptor_memory_s1_begins_xfer = ~d1_reasons_to_wait & ((pb_cpu_to_io_m1_qualified_request_descriptor_memory_s1 | pb_dma_to_descriptor_memory_m1_qualified_request_descriptor_memory_s1));
  //assign descriptor_memory_s1_readdata_from_sa = descriptor_memory_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign descriptor_memory_s1_readdata_from_sa = descriptor_memory_s1_readdata;

  assign pb_cpu_to_io_m1_requests_descriptor_memory_s1 = ({pb_cpu_to_io_m1_address_to_slave[22 : 13] , 13'b0} == 23'h2000) & pb_cpu_to_io_m1_chipselect;
  //descriptor_memory_s1_arb_share_counter set values, which is an e_mux
  assign descriptor_memory_s1_arb_share_set_values = (pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1)? 8 :
    (pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1)? 8 :
    1;

  //descriptor_memory_s1_non_bursting_master_requests mux, which is an e_mux
  assign descriptor_memory_s1_non_bursting_master_requests = pb_cpu_to_io_m1_requests_descriptor_memory_s1 |
    pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1 |
    pb_cpu_to_io_m1_requests_descriptor_memory_s1 |
    pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1;

  //descriptor_memory_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign descriptor_memory_s1_any_bursting_master_saved_grant = 0;

  //descriptor_memory_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign descriptor_memory_s1_arb_share_counter_next_value = descriptor_memory_s1_firsttransfer ? (descriptor_memory_s1_arb_share_set_values - 1) : |descriptor_memory_s1_arb_share_counter ? (descriptor_memory_s1_arb_share_counter - 1) : 0;

  //descriptor_memory_s1_allgrants all slave grants, which is an e_mux
  assign descriptor_memory_s1_allgrants = (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector);

  //descriptor_memory_s1_end_xfer assignment, which is an e_assign
  assign descriptor_memory_s1_end_xfer = ~(descriptor_memory_s1_waits_for_read | descriptor_memory_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_descriptor_memory_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_descriptor_memory_s1 = descriptor_memory_s1_end_xfer & (~descriptor_memory_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //descriptor_memory_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign descriptor_memory_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_descriptor_memory_s1 & descriptor_memory_s1_allgrants) | (end_xfer_arb_share_counter_term_descriptor_memory_s1 & ~descriptor_memory_s1_non_bursting_master_requests);

  //descriptor_memory_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_arb_share_counter <= 0;
      else if (descriptor_memory_s1_arb_counter_enable)
          descriptor_memory_s1_arb_share_counter <= descriptor_memory_s1_arb_share_counter_next_value;
    end


  //descriptor_memory_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_slavearbiterlockenable <= 0;
      else if ((|descriptor_memory_s1_master_qreq_vector & end_xfer_arb_share_counter_term_descriptor_memory_s1) | (end_xfer_arb_share_counter_term_descriptor_memory_s1 & ~descriptor_memory_s1_non_bursting_master_requests))
          descriptor_memory_s1_slavearbiterlockenable <= |descriptor_memory_s1_arb_share_counter_next_value;
    end


  //pb_cpu_to_io/m1 descriptor_memory/s1 arbiterlock, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock = descriptor_memory_s1_slavearbiterlockenable & pb_cpu_to_io_m1_continuerequest;

  //descriptor_memory_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign descriptor_memory_s1_slavearbiterlockenable2 = |descriptor_memory_s1_arb_share_counter_next_value;

  //pb_cpu_to_io/m1 descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock2 = descriptor_memory_s1_slavearbiterlockenable2 & pb_cpu_to_io_m1_continuerequest;

  //pb_dma_to_descriptor_memory/m1 descriptor_memory/s1 arbiterlock, which is an e_assign
  assign pb_dma_to_descriptor_memory_m1_arbiterlock = descriptor_memory_s1_slavearbiterlockenable & pb_dma_to_descriptor_memory_m1_continuerequest;

  //pb_dma_to_descriptor_memory/m1 descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign pb_dma_to_descriptor_memory_m1_arbiterlock2 = descriptor_memory_s1_slavearbiterlockenable2 & pb_dma_to_descriptor_memory_m1_continuerequest;

  //pb_dma_to_descriptor_memory/m1 granted descriptor_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_pb_dma_to_descriptor_memory_m1_granted_slave_descriptor_memory_s1 <= 0;
      else 
        last_cycle_pb_dma_to_descriptor_memory_m1_granted_slave_descriptor_memory_s1 <= pb_dma_to_descriptor_memory_m1_saved_grant_descriptor_memory_s1 ? 1 : (descriptor_memory_s1_arbitration_holdoff_internal | ~pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1) ? 0 : last_cycle_pb_dma_to_descriptor_memory_m1_granted_slave_descriptor_memory_s1;
    end


  //pb_dma_to_descriptor_memory_m1_continuerequest continued request, which is an e_mux
  assign pb_dma_to_descriptor_memory_m1_continuerequest = last_cycle_pb_dma_to_descriptor_memory_m1_granted_slave_descriptor_memory_s1 & pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1;

  //descriptor_memory_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign descriptor_memory_s1_any_continuerequest = pb_dma_to_descriptor_memory_m1_continuerequest |
    pb_cpu_to_io_m1_continuerequest;

  assign pb_cpu_to_io_m1_qualified_request_descriptor_memory_s1 = pb_cpu_to_io_m1_requests_descriptor_memory_s1 & ~(((pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ((1 < pb_cpu_to_io_m1_latency_counter))) | pb_dma_to_descriptor_memory_m1_arbiterlock);
  //pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1_shift_register_in = pb_cpu_to_io_m1_granted_descriptor_memory_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ~descriptor_memory_s1_waits_for_read;

  //shift register p1 pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1_shift_register = {pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1_shift_register, pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1_shift_register_in};

  //pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1_shift_register <= 0;
      else 
        pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1_shift_register <= p1_pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1_shift_register;
    end


  //local readdatavalid pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1, which is an e_mux
  assign pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1 = pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1_shift_register;

  //descriptor_memory_s1_writedata mux, which is an e_mux
  assign descriptor_memory_s1_writedata = (pb_cpu_to_io_m1_granted_descriptor_memory_s1)? pb_cpu_to_io_m1_writedata :
    pb_dma_to_descriptor_memory_m1_writedata;

  //mux descriptor_memory_s1_clken, which is an e_mux
  assign descriptor_memory_s1_clken = 1'b1;

  assign pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1 = ({pb_dma_to_descriptor_memory_m1_address_to_slave[13] , 13'b0} == 14'h2000) & pb_dma_to_descriptor_memory_m1_chipselect;
  //pb_cpu_to_io/m1 granted descriptor_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_pb_cpu_to_io_m1_granted_slave_descriptor_memory_s1 <= 0;
      else 
        last_cycle_pb_cpu_to_io_m1_granted_slave_descriptor_memory_s1 <= pb_cpu_to_io_m1_saved_grant_descriptor_memory_s1 ? 1 : (descriptor_memory_s1_arbitration_holdoff_internal | ~pb_cpu_to_io_m1_requests_descriptor_memory_s1) ? 0 : last_cycle_pb_cpu_to_io_m1_granted_slave_descriptor_memory_s1;
    end


  //pb_cpu_to_io_m1_continuerequest continued request, which is an e_mux
  assign pb_cpu_to_io_m1_continuerequest = last_cycle_pb_cpu_to_io_m1_granted_slave_descriptor_memory_s1 & pb_cpu_to_io_m1_requests_descriptor_memory_s1;

  assign pb_dma_to_descriptor_memory_m1_qualified_request_descriptor_memory_s1 = pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1 & ~(pb_cpu_to_io_m1_arbiterlock);
  //pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1_shift_register_in = pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1 & (pb_dma_to_descriptor_memory_m1_read & pb_dma_to_descriptor_memory_m1_chipselect) & ~descriptor_memory_s1_waits_for_read;

  //shift register p1 pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1_shift_register = {pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1_shift_register, pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1_shift_register_in};

  //pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1_shift_register <= 0;
      else 
        pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1_shift_register <= p1_pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1_shift_register;
    end


  //local readdatavalid pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1, which is an e_mux
  assign pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1 = pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1_shift_register;

  //allow new arb cycle for descriptor_memory/s1, which is an e_assign
  assign descriptor_memory_s1_allow_new_arb_cycle = ~pb_cpu_to_io_m1_arbiterlock & ~pb_dma_to_descriptor_memory_m1_arbiterlock;

  //pb_dma_to_descriptor_memory/m1 assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  assign descriptor_memory_s1_master_qreq_vector[0] = pb_dma_to_descriptor_memory_m1_qualified_request_descriptor_memory_s1;

  //pb_dma_to_descriptor_memory/m1 grant descriptor_memory/s1, which is an e_assign
  assign pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1 = descriptor_memory_s1_grant_vector[0];

  //pb_dma_to_descriptor_memory/m1 saved-grant descriptor_memory/s1, which is an e_assign
  assign pb_dma_to_descriptor_memory_m1_saved_grant_descriptor_memory_s1 = descriptor_memory_s1_arb_winner[0] && pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1;

  //pb_cpu_to_io/m1 assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  assign descriptor_memory_s1_master_qreq_vector[1] = pb_cpu_to_io_m1_qualified_request_descriptor_memory_s1;

  //pb_cpu_to_io/m1 grant descriptor_memory/s1, which is an e_assign
  assign pb_cpu_to_io_m1_granted_descriptor_memory_s1 = descriptor_memory_s1_grant_vector[1];

  //pb_cpu_to_io/m1 saved-grant descriptor_memory/s1, which is an e_assign
  assign pb_cpu_to_io_m1_saved_grant_descriptor_memory_s1 = descriptor_memory_s1_arb_winner[1] && pb_cpu_to_io_m1_requests_descriptor_memory_s1;

  //descriptor_memory/s1 chosen-master double-vector, which is an e_assign
  assign descriptor_memory_s1_chosen_master_double_vector = {descriptor_memory_s1_master_qreq_vector, descriptor_memory_s1_master_qreq_vector} & ({~descriptor_memory_s1_master_qreq_vector, ~descriptor_memory_s1_master_qreq_vector} + descriptor_memory_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign descriptor_memory_s1_arb_winner = (descriptor_memory_s1_allow_new_arb_cycle & | descriptor_memory_s1_grant_vector) ? descriptor_memory_s1_grant_vector : descriptor_memory_s1_saved_chosen_master_vector;

  //saved descriptor_memory_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_saved_chosen_master_vector <= 0;
      else if (descriptor_memory_s1_allow_new_arb_cycle)
          descriptor_memory_s1_saved_chosen_master_vector <= |descriptor_memory_s1_grant_vector ? descriptor_memory_s1_grant_vector : descriptor_memory_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign descriptor_memory_s1_grant_vector = {(descriptor_memory_s1_chosen_master_double_vector[1] | descriptor_memory_s1_chosen_master_double_vector[3]),
    (descriptor_memory_s1_chosen_master_double_vector[0] | descriptor_memory_s1_chosen_master_double_vector[2])};

  //descriptor_memory/s1 chosen master rotated left, which is an e_assign
  assign descriptor_memory_s1_chosen_master_rot_left = (descriptor_memory_s1_arb_winner << 1) ? (descriptor_memory_s1_arb_winner << 1) : 1;

  //descriptor_memory/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_arb_addend <= 1;
      else if (|descriptor_memory_s1_grant_vector)
          descriptor_memory_s1_arb_addend <= descriptor_memory_s1_end_xfer? descriptor_memory_s1_chosen_master_rot_left : descriptor_memory_s1_grant_vector;
    end


  //~descriptor_memory_s1_reset assignment, which is an e_assign
  assign descriptor_memory_s1_reset = ~reset_n;

  assign descriptor_memory_s1_chipselect = pb_cpu_to_io_m1_granted_descriptor_memory_s1 | pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1;
  //descriptor_memory_s1_firsttransfer first transaction, which is an e_assign
  assign descriptor_memory_s1_firsttransfer = descriptor_memory_s1_begins_xfer ? descriptor_memory_s1_unreg_firsttransfer : descriptor_memory_s1_reg_firsttransfer;

  //descriptor_memory_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign descriptor_memory_s1_unreg_firsttransfer = ~(descriptor_memory_s1_slavearbiterlockenable & descriptor_memory_s1_any_continuerequest);

  //descriptor_memory_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_reg_firsttransfer <= 1'b1;
      else if (descriptor_memory_s1_begins_xfer)
          descriptor_memory_s1_reg_firsttransfer <= descriptor_memory_s1_unreg_firsttransfer;
    end


  //descriptor_memory_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign descriptor_memory_s1_beginbursttransfer_internal = descriptor_memory_s1_begins_xfer;

  //descriptor_memory_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign descriptor_memory_s1_arbitration_holdoff_internal = descriptor_memory_s1_begins_xfer & descriptor_memory_s1_firsttransfer;

  //descriptor_memory_s1_write assignment, which is an e_mux
  assign descriptor_memory_s1_write = (pb_cpu_to_io_m1_granted_descriptor_memory_s1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect)) | (pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1 & (pb_dma_to_descriptor_memory_m1_write & pb_dma_to_descriptor_memory_m1_chipselect));

  assign shifted_address_to_descriptor_memory_s1_from_pb_cpu_to_io_m1 = pb_cpu_to_io_m1_address_to_slave;
  //descriptor_memory_s1_address mux, which is an e_mux
  assign descriptor_memory_s1_address = (pb_cpu_to_io_m1_granted_descriptor_memory_s1)? (shifted_address_to_descriptor_memory_s1_from_pb_cpu_to_io_m1 >> 2) :
    (shifted_address_to_descriptor_memory_s1_from_pb_dma_to_descriptor_memory_m1 >> 2);

  assign shifted_address_to_descriptor_memory_s1_from_pb_dma_to_descriptor_memory_m1 = pb_dma_to_descriptor_memory_m1_address_to_slave;
  //d1_descriptor_memory_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_descriptor_memory_s1_end_xfer <= 1;
      else 
        d1_descriptor_memory_s1_end_xfer <= descriptor_memory_s1_end_xfer;
    end


  //descriptor_memory_s1_waits_for_read in a cycle, which is an e_mux
  assign descriptor_memory_s1_waits_for_read = descriptor_memory_s1_in_a_read_cycle & 0;

  //descriptor_memory_s1_in_a_read_cycle assignment, which is an e_assign
  assign descriptor_memory_s1_in_a_read_cycle = (pb_cpu_to_io_m1_granted_descriptor_memory_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)) | (pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1 & (pb_dma_to_descriptor_memory_m1_read & pb_dma_to_descriptor_memory_m1_chipselect));

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = descriptor_memory_s1_in_a_read_cycle;

  //descriptor_memory_s1_waits_for_write in a cycle, which is an e_mux
  assign descriptor_memory_s1_waits_for_write = descriptor_memory_s1_in_a_write_cycle & 0;

  //descriptor_memory_s1_in_a_write_cycle assignment, which is an e_assign
  assign descriptor_memory_s1_in_a_write_cycle = (pb_cpu_to_io_m1_granted_descriptor_memory_s1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect)) | (pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1 & (pb_dma_to_descriptor_memory_m1_write & pb_dma_to_descriptor_memory_m1_chipselect));

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = descriptor_memory_s1_in_a_write_cycle;

  assign wait_for_descriptor_memory_s1_counter = 0;
  //descriptor_memory_s1_byteenable byte enable port mux, which is an e_mux
  assign descriptor_memory_s1_byteenable = (pb_cpu_to_io_m1_granted_descriptor_memory_s1)? pb_cpu_to_io_m1_byteenable :
    (pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1)? pb_dma_to_descriptor_memory_m1_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //descriptor_memory/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pb_cpu_to_io/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_io_m1_requests_descriptor_memory_s1 && (pb_cpu_to_io_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pb_cpu_to_io/m1 drove 0 on its 'burstcount' port while accessing slave descriptor_memory/s1", $time);
          $stop;
        end
    end


  //pb_dma_to_descriptor_memory/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1 && (pb_dma_to_descriptor_memory_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pb_dma_to_descriptor_memory/m1 drove 0 on its 'burstcount' port while accessing slave descriptor_memory/s1", $time);
          $stop;
        end
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_io_m1_granted_descriptor_memory_s1 + pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_io_m1_saved_grant_descriptor_memory_s1 + pb_dma_to_descriptor_memory_m1_saved_grant_descriptor_memory_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module dipsw_pio_s1_arbitrator (
                                 // inputs:
                                  clk,
                                  dipsw_pio_s1_irq,
                                  dipsw_pio_s1_readdata,
                                  pb_cpu_to_io_m1_address_to_slave,
                                  pb_cpu_to_io_m1_burstcount,
                                  pb_cpu_to_io_m1_byteenable,
                                  pb_cpu_to_io_m1_chipselect,
                                  pb_cpu_to_io_m1_latency_counter,
                                  pb_cpu_to_io_m1_read,
                                  pb_cpu_to_io_m1_write,
                                  pb_cpu_to_io_m1_writedata,
                                  reset_n,

                                 // outputs:
                                  d1_dipsw_pio_s1_end_xfer,
                                  dipsw_pio_s1_address,
                                  dipsw_pio_s1_chipselect,
                                  dipsw_pio_s1_irq_from_sa,
                                  dipsw_pio_s1_readdata_from_sa,
                                  dipsw_pio_s1_reset_n,
                                  dipsw_pio_s1_write_n,
                                  dipsw_pio_s1_writedata,
                                  pb_cpu_to_io_m1_granted_dipsw_pio_s1,
                                  pb_cpu_to_io_m1_qualified_request_dipsw_pio_s1,
                                  pb_cpu_to_io_m1_read_data_valid_dipsw_pio_s1,
                                  pb_cpu_to_io_m1_requests_dipsw_pio_s1
                               )
;

  output           d1_dipsw_pio_s1_end_xfer;
  output  [  1: 0] dipsw_pio_s1_address;
  output           dipsw_pio_s1_chipselect;
  output           dipsw_pio_s1_irq_from_sa;
  output  [  7: 0] dipsw_pio_s1_readdata_from_sa;
  output           dipsw_pio_s1_reset_n;
  output           dipsw_pio_s1_write_n;
  output  [  7: 0] dipsw_pio_s1_writedata;
  output           pb_cpu_to_io_m1_granted_dipsw_pio_s1;
  output           pb_cpu_to_io_m1_qualified_request_dipsw_pio_s1;
  output           pb_cpu_to_io_m1_read_data_valid_dipsw_pio_s1;
  output           pb_cpu_to_io_m1_requests_dipsw_pio_s1;
  input            clk;
  input            dipsw_pio_s1_irq;
  input   [  7: 0] dipsw_pio_s1_readdata;
  input   [ 22: 0] pb_cpu_to_io_m1_address_to_slave;
  input            pb_cpu_to_io_m1_burstcount;
  input   [  3: 0] pb_cpu_to_io_m1_byteenable;
  input            pb_cpu_to_io_m1_chipselect;
  input            pb_cpu_to_io_m1_latency_counter;
  input            pb_cpu_to_io_m1_read;
  input            pb_cpu_to_io_m1_write;
  input   [ 31: 0] pb_cpu_to_io_m1_writedata;
  input            reset_n;

  reg              d1_dipsw_pio_s1_end_xfer;
  reg              d1_reasons_to_wait;
  wire    [  1: 0] dipsw_pio_s1_address;
  wire             dipsw_pio_s1_allgrants;
  wire             dipsw_pio_s1_allow_new_arb_cycle;
  wire             dipsw_pio_s1_any_bursting_master_saved_grant;
  wire             dipsw_pio_s1_any_continuerequest;
  wire             dipsw_pio_s1_arb_counter_enable;
  reg              dipsw_pio_s1_arb_share_counter;
  wire             dipsw_pio_s1_arb_share_counter_next_value;
  wire             dipsw_pio_s1_arb_share_set_values;
  wire             dipsw_pio_s1_beginbursttransfer_internal;
  wire             dipsw_pio_s1_begins_xfer;
  wire             dipsw_pio_s1_chipselect;
  wire             dipsw_pio_s1_end_xfer;
  wire             dipsw_pio_s1_firsttransfer;
  wire             dipsw_pio_s1_grant_vector;
  wire             dipsw_pio_s1_in_a_read_cycle;
  wire             dipsw_pio_s1_in_a_write_cycle;
  wire             dipsw_pio_s1_irq_from_sa;
  wire             dipsw_pio_s1_master_qreq_vector;
  wire             dipsw_pio_s1_non_bursting_master_requests;
  wire             dipsw_pio_s1_pretend_byte_enable;
  wire    [  7: 0] dipsw_pio_s1_readdata_from_sa;
  reg              dipsw_pio_s1_reg_firsttransfer;
  wire             dipsw_pio_s1_reset_n;
  reg              dipsw_pio_s1_slavearbiterlockenable;
  wire             dipsw_pio_s1_slavearbiterlockenable2;
  wire             dipsw_pio_s1_unreg_firsttransfer;
  wire             dipsw_pio_s1_waits_for_read;
  wire             dipsw_pio_s1_waits_for_write;
  wire             dipsw_pio_s1_write_n;
  wire    [  7: 0] dipsw_pio_s1_writedata;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_dipsw_pio_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             pb_cpu_to_io_m1_arbiterlock;
  wire             pb_cpu_to_io_m1_arbiterlock2;
  wire             pb_cpu_to_io_m1_continuerequest;
  wire             pb_cpu_to_io_m1_granted_dipsw_pio_s1;
  wire             pb_cpu_to_io_m1_qualified_request_dipsw_pio_s1;
  wire             pb_cpu_to_io_m1_read_data_valid_dipsw_pio_s1;
  wire             pb_cpu_to_io_m1_requests_dipsw_pio_s1;
  wire             pb_cpu_to_io_m1_saved_grant_dipsw_pio_s1;
  wire    [ 22: 0] shifted_address_to_dipsw_pio_s1_from_pb_cpu_to_io_m1;
  wire             wait_for_dipsw_pio_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~dipsw_pio_s1_end_xfer;
    end


  assign dipsw_pio_s1_begins_xfer = ~d1_reasons_to_wait & ((pb_cpu_to_io_m1_qualified_request_dipsw_pio_s1));
  //assign dipsw_pio_s1_readdata_from_sa = dipsw_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign dipsw_pio_s1_readdata_from_sa = dipsw_pio_s1_readdata;

  assign pb_cpu_to_io_m1_requests_dipsw_pio_s1 = ({pb_cpu_to_io_m1_address_to_slave[22 : 4] , 4'b0} == 23'h4ce0) & pb_cpu_to_io_m1_chipselect;
  //dipsw_pio_s1_arb_share_counter set values, which is an e_mux
  assign dipsw_pio_s1_arb_share_set_values = 1;

  //dipsw_pio_s1_non_bursting_master_requests mux, which is an e_mux
  assign dipsw_pio_s1_non_bursting_master_requests = pb_cpu_to_io_m1_requests_dipsw_pio_s1;

  //dipsw_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign dipsw_pio_s1_any_bursting_master_saved_grant = 0;

  //dipsw_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign dipsw_pio_s1_arb_share_counter_next_value = dipsw_pio_s1_firsttransfer ? (dipsw_pio_s1_arb_share_set_values - 1) : |dipsw_pio_s1_arb_share_counter ? (dipsw_pio_s1_arb_share_counter - 1) : 0;

  //dipsw_pio_s1_allgrants all slave grants, which is an e_mux
  assign dipsw_pio_s1_allgrants = |dipsw_pio_s1_grant_vector;

  //dipsw_pio_s1_end_xfer assignment, which is an e_assign
  assign dipsw_pio_s1_end_xfer = ~(dipsw_pio_s1_waits_for_read | dipsw_pio_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_dipsw_pio_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_dipsw_pio_s1 = dipsw_pio_s1_end_xfer & (~dipsw_pio_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //dipsw_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign dipsw_pio_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_dipsw_pio_s1 & dipsw_pio_s1_allgrants) | (end_xfer_arb_share_counter_term_dipsw_pio_s1 & ~dipsw_pio_s1_non_bursting_master_requests);

  //dipsw_pio_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dipsw_pio_s1_arb_share_counter <= 0;
      else if (dipsw_pio_s1_arb_counter_enable)
          dipsw_pio_s1_arb_share_counter <= dipsw_pio_s1_arb_share_counter_next_value;
    end


  //dipsw_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dipsw_pio_s1_slavearbiterlockenable <= 0;
      else if ((|dipsw_pio_s1_master_qreq_vector & end_xfer_arb_share_counter_term_dipsw_pio_s1) | (end_xfer_arb_share_counter_term_dipsw_pio_s1 & ~dipsw_pio_s1_non_bursting_master_requests))
          dipsw_pio_s1_slavearbiterlockenable <= |dipsw_pio_s1_arb_share_counter_next_value;
    end


  //pb_cpu_to_io/m1 dipsw_pio/s1 arbiterlock, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock = dipsw_pio_s1_slavearbiterlockenable & pb_cpu_to_io_m1_continuerequest;

  //dipsw_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign dipsw_pio_s1_slavearbiterlockenable2 = |dipsw_pio_s1_arb_share_counter_next_value;

  //pb_cpu_to_io/m1 dipsw_pio/s1 arbiterlock2, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock2 = dipsw_pio_s1_slavearbiterlockenable2 & pb_cpu_to_io_m1_continuerequest;

  //dipsw_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign dipsw_pio_s1_any_continuerequest = 1;

  //pb_cpu_to_io_m1_continuerequest continued request, which is an e_assign
  assign pb_cpu_to_io_m1_continuerequest = 1;

  assign pb_cpu_to_io_m1_qualified_request_dipsw_pio_s1 = pb_cpu_to_io_m1_requests_dipsw_pio_s1 & ~(((pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ((pb_cpu_to_io_m1_latency_counter != 0))));
  //local readdatavalid pb_cpu_to_io_m1_read_data_valid_dipsw_pio_s1, which is an e_mux
  assign pb_cpu_to_io_m1_read_data_valid_dipsw_pio_s1 = pb_cpu_to_io_m1_granted_dipsw_pio_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ~dipsw_pio_s1_waits_for_read;

  //dipsw_pio_s1_writedata mux, which is an e_mux
  assign dipsw_pio_s1_writedata = pb_cpu_to_io_m1_writedata;

  //master is always granted when requested
  assign pb_cpu_to_io_m1_granted_dipsw_pio_s1 = pb_cpu_to_io_m1_qualified_request_dipsw_pio_s1;

  //pb_cpu_to_io/m1 saved-grant dipsw_pio/s1, which is an e_assign
  assign pb_cpu_to_io_m1_saved_grant_dipsw_pio_s1 = pb_cpu_to_io_m1_requests_dipsw_pio_s1;

  //allow new arb cycle for dipsw_pio/s1, which is an e_assign
  assign dipsw_pio_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign dipsw_pio_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign dipsw_pio_s1_master_qreq_vector = 1;

  //dipsw_pio_s1_reset_n assignment, which is an e_assign
  assign dipsw_pio_s1_reset_n = reset_n;

  assign dipsw_pio_s1_chipselect = pb_cpu_to_io_m1_granted_dipsw_pio_s1;
  //dipsw_pio_s1_firsttransfer first transaction, which is an e_assign
  assign dipsw_pio_s1_firsttransfer = dipsw_pio_s1_begins_xfer ? dipsw_pio_s1_unreg_firsttransfer : dipsw_pio_s1_reg_firsttransfer;

  //dipsw_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign dipsw_pio_s1_unreg_firsttransfer = ~(dipsw_pio_s1_slavearbiterlockenable & dipsw_pio_s1_any_continuerequest);

  //dipsw_pio_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dipsw_pio_s1_reg_firsttransfer <= 1'b1;
      else if (dipsw_pio_s1_begins_xfer)
          dipsw_pio_s1_reg_firsttransfer <= dipsw_pio_s1_unreg_firsttransfer;
    end


  //dipsw_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign dipsw_pio_s1_beginbursttransfer_internal = dipsw_pio_s1_begins_xfer;

  //~dipsw_pio_s1_write_n assignment, which is an e_mux
  assign dipsw_pio_s1_write_n = ~(((pb_cpu_to_io_m1_granted_dipsw_pio_s1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect))) & dipsw_pio_s1_pretend_byte_enable);

  assign shifted_address_to_dipsw_pio_s1_from_pb_cpu_to_io_m1 = pb_cpu_to_io_m1_address_to_slave;
  //dipsw_pio_s1_address mux, which is an e_mux
  assign dipsw_pio_s1_address = shifted_address_to_dipsw_pio_s1_from_pb_cpu_to_io_m1 >> 2;

  //d1_dipsw_pio_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_dipsw_pio_s1_end_xfer <= 1;
      else 
        d1_dipsw_pio_s1_end_xfer <= dipsw_pio_s1_end_xfer;
    end


  //dipsw_pio_s1_waits_for_read in a cycle, which is an e_mux
  assign dipsw_pio_s1_waits_for_read = dipsw_pio_s1_in_a_read_cycle & dipsw_pio_s1_begins_xfer;

  //dipsw_pio_s1_in_a_read_cycle assignment, which is an e_assign
  assign dipsw_pio_s1_in_a_read_cycle = pb_cpu_to_io_m1_granted_dipsw_pio_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = dipsw_pio_s1_in_a_read_cycle;

  //dipsw_pio_s1_waits_for_write in a cycle, which is an e_mux
  assign dipsw_pio_s1_waits_for_write = dipsw_pio_s1_in_a_write_cycle & 0;

  //dipsw_pio_s1_in_a_write_cycle assignment, which is an e_assign
  assign dipsw_pio_s1_in_a_write_cycle = pb_cpu_to_io_m1_granted_dipsw_pio_s1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = dipsw_pio_s1_in_a_write_cycle;

  assign wait_for_dipsw_pio_s1_counter = 0;
  //dipsw_pio_s1_pretend_byte_enable byte enable port mux, which is an e_mux
  assign dipsw_pio_s1_pretend_byte_enable = (pb_cpu_to_io_m1_granted_dipsw_pio_s1)? pb_cpu_to_io_m1_byteenable :
    -1;

  //assign dipsw_pio_s1_irq_from_sa = dipsw_pio_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign dipsw_pio_s1_irq_from_sa = dipsw_pio_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //dipsw_pio/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pb_cpu_to_io/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_io_m1_requests_dipsw_pio_s1 && (pb_cpu_to_io_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pb_cpu_to_io/m1 drove 0 on its 'burstcount' port while accessing slave dipsw_pio/s1", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_avalon_jtag_slave_arbitrator (
                                                // inputs:
                                                 clk,
                                                 jtag_uart_avalon_jtag_slave_dataavailable,
                                                 jtag_uart_avalon_jtag_slave_irq,
                                                 jtag_uart_avalon_jtag_slave_readdata,
                                                 jtag_uart_avalon_jtag_slave_readyfordata,
                                                 jtag_uart_avalon_jtag_slave_waitrequest,
                                                 pb_cpu_to_io_m1_address_to_slave,
                                                 pb_cpu_to_io_m1_burstcount,
                                                 pb_cpu_to_io_m1_chipselect,
                                                 pb_cpu_to_io_m1_latency_counter,
                                                 pb_cpu_to_io_m1_read,
                                                 pb_cpu_to_io_m1_write,
                                                 pb_cpu_to_io_m1_writedata,
                                                 reset_n,

                                                // outputs:
                                                 d1_jtag_uart_avalon_jtag_slave_end_xfer,
                                                 jtag_uart_avalon_jtag_slave_address,
                                                 jtag_uart_avalon_jtag_slave_chipselect,
                                                 jtag_uart_avalon_jtag_slave_dataavailable_from_sa,
                                                 jtag_uart_avalon_jtag_slave_irq_from_sa,
                                                 jtag_uart_avalon_jtag_slave_read_n,
                                                 jtag_uart_avalon_jtag_slave_readdata_from_sa,
                                                 jtag_uart_avalon_jtag_slave_readyfordata_from_sa,
                                                 jtag_uart_avalon_jtag_slave_reset_n,
                                                 jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
                                                 jtag_uart_avalon_jtag_slave_write_n,
                                                 jtag_uart_avalon_jtag_slave_writedata,
                                                 pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave,
                                                 pb_cpu_to_io_m1_qualified_request_jtag_uart_avalon_jtag_slave,
                                                 pb_cpu_to_io_m1_read_data_valid_jtag_uart_avalon_jtag_slave,
                                                 pb_cpu_to_io_m1_requests_jtag_uart_avalon_jtag_slave
                                              )
;

  output           d1_jtag_uart_avalon_jtag_slave_end_xfer;
  output           jtag_uart_avalon_jtag_slave_address;
  output           jtag_uart_avalon_jtag_slave_chipselect;
  output           jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  output           jtag_uart_avalon_jtag_slave_irq_from_sa;
  output           jtag_uart_avalon_jtag_slave_read_n;
  output  [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  output           jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  output           jtag_uart_avalon_jtag_slave_reset_n;
  output           jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  output           jtag_uart_avalon_jtag_slave_write_n;
  output  [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  output           pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave;
  output           pb_cpu_to_io_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  output           pb_cpu_to_io_m1_read_data_valid_jtag_uart_avalon_jtag_slave;
  output           pb_cpu_to_io_m1_requests_jtag_uart_avalon_jtag_slave;
  input            clk;
  input            jtag_uart_avalon_jtag_slave_dataavailable;
  input            jtag_uart_avalon_jtag_slave_irq;
  input   [ 31: 0] jtag_uart_avalon_jtag_slave_readdata;
  input            jtag_uart_avalon_jtag_slave_readyfordata;
  input            jtag_uart_avalon_jtag_slave_waitrequest;
  input   [ 22: 0] pb_cpu_to_io_m1_address_to_slave;
  input            pb_cpu_to_io_m1_burstcount;
  input            pb_cpu_to_io_m1_chipselect;
  input            pb_cpu_to_io_m1_latency_counter;
  input            pb_cpu_to_io_m1_read;
  input            pb_cpu_to_io_m1_write;
  input   [ 31: 0] pb_cpu_to_io_m1_writedata;
  input            reset_n;

  reg              d1_jtag_uart_avalon_jtag_slave_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             jtag_uart_avalon_jtag_slave_address;
  wire             jtag_uart_avalon_jtag_slave_allgrants;
  wire             jtag_uart_avalon_jtag_slave_allow_new_arb_cycle;
  wire             jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant;
  wire             jtag_uart_avalon_jtag_slave_any_continuerequest;
  wire             jtag_uart_avalon_jtag_slave_arb_counter_enable;
  reg              jtag_uart_avalon_jtag_slave_arb_share_counter;
  wire             jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
  wire             jtag_uart_avalon_jtag_slave_arb_share_set_values;
  wire             jtag_uart_avalon_jtag_slave_beginbursttransfer_internal;
  wire             jtag_uart_avalon_jtag_slave_begins_xfer;
  wire             jtag_uart_avalon_jtag_slave_chipselect;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_end_xfer;
  wire             jtag_uart_avalon_jtag_slave_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_grant_vector;
  wire             jtag_uart_avalon_jtag_slave_in_a_read_cycle;
  wire             jtag_uart_avalon_jtag_slave_in_a_write_cycle;
  wire             jtag_uart_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_avalon_jtag_slave_master_qreq_vector;
  wire             jtag_uart_avalon_jtag_slave_non_bursting_master_requests;
  wire             jtag_uart_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  reg              jtag_uart_avalon_jtag_slave_reg_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_reset_n;
  reg              jtag_uart_avalon_jtag_slave_slavearbiterlockenable;
  wire             jtag_uart_avalon_jtag_slave_slavearbiterlockenable2;
  wire             jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_avalon_jtag_slave_waits_for_read;
  wire             jtag_uart_avalon_jtag_slave_waits_for_write;
  wire             jtag_uart_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  wire             pb_cpu_to_io_m1_arbiterlock;
  wire             pb_cpu_to_io_m1_arbiterlock2;
  wire             pb_cpu_to_io_m1_continuerequest;
  wire             pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave;
  wire             pb_cpu_to_io_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  wire             pb_cpu_to_io_m1_read_data_valid_jtag_uart_avalon_jtag_slave;
  wire             pb_cpu_to_io_m1_requests_jtag_uart_avalon_jtag_slave;
  wire             pb_cpu_to_io_m1_saved_grant_jtag_uart_avalon_jtag_slave;
  wire    [ 22: 0] shifted_address_to_jtag_uart_avalon_jtag_slave_from_pb_cpu_to_io_m1;
  wire             wait_for_jtag_uart_avalon_jtag_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~jtag_uart_avalon_jtag_slave_end_xfer;
    end


  assign jtag_uart_avalon_jtag_slave_begins_xfer = ~d1_reasons_to_wait & ((pb_cpu_to_io_m1_qualified_request_jtag_uart_avalon_jtag_slave));
  //assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata;

  assign pb_cpu_to_io_m1_requests_jtag_uart_avalon_jtag_slave = ({pb_cpu_to_io_m1_address_to_slave[22 : 3] , 3'b0} == 23'h4d50) & pb_cpu_to_io_m1_chipselect;
  //assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable;

  //assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata;

  //assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest;

  //jtag_uart_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_arb_share_set_values = 1;

  //jtag_uart_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_non_bursting_master_requests = pb_cpu_to_io_m1_requests_jtag_uart_avalon_jtag_slave;

  //jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant = 0;

  //jtag_uart_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_arb_share_counter_next_value = jtag_uart_avalon_jtag_slave_firsttransfer ? (jtag_uart_avalon_jtag_slave_arb_share_set_values - 1) : |jtag_uart_avalon_jtag_slave_arb_share_counter ? (jtag_uart_avalon_jtag_slave_arb_share_counter - 1) : 0;

  //jtag_uart_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_allgrants = |jtag_uart_avalon_jtag_slave_grant_vector;

  //jtag_uart_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_end_xfer = ~(jtag_uart_avalon_jtag_slave_waits_for_read | jtag_uart_avalon_jtag_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave = jtag_uart_avalon_jtag_slave_end_xfer & (~jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //jtag_uart_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & jtag_uart_avalon_jtag_slave_allgrants) | (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & ~jtag_uart_avalon_jtag_slave_non_bursting_master_requests);

  //jtag_uart_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_arb_share_counter <= 0;
      else if (jtag_uart_avalon_jtag_slave_arb_counter_enable)
          jtag_uart_avalon_jtag_slave_arb_share_counter <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //jtag_uart_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= 0;
      else if ((|jtag_uart_avalon_jtag_slave_master_qreq_vector & end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave) | (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & ~jtag_uart_avalon_jtag_slave_non_bursting_master_requests))
          jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= |jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //pb_cpu_to_io/m1 jtag_uart/avalon_jtag_slave arbiterlock, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock = jtag_uart_avalon_jtag_slave_slavearbiterlockenable & pb_cpu_to_io_m1_continuerequest;

  //jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 = |jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;

  //pb_cpu_to_io/m1 jtag_uart/avalon_jtag_slave arbiterlock2, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock2 = jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 & pb_cpu_to_io_m1_continuerequest;

  //jtag_uart_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_any_continuerequest = 1;

  //pb_cpu_to_io_m1_continuerequest continued request, which is an e_assign
  assign pb_cpu_to_io_m1_continuerequest = 1;

  assign pb_cpu_to_io_m1_qualified_request_jtag_uart_avalon_jtag_slave = pb_cpu_to_io_m1_requests_jtag_uart_avalon_jtag_slave & ~(((pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ((pb_cpu_to_io_m1_latency_counter != 0))));
  //local readdatavalid pb_cpu_to_io_m1_read_data_valid_jtag_uart_avalon_jtag_slave, which is an e_mux
  assign pb_cpu_to_io_m1_read_data_valid_jtag_uart_avalon_jtag_slave = pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ~jtag_uart_avalon_jtag_slave_waits_for_read;

  //jtag_uart_avalon_jtag_slave_writedata mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_writedata = pb_cpu_to_io_m1_writedata;

  //master is always granted when requested
  assign pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave = pb_cpu_to_io_m1_qualified_request_jtag_uart_avalon_jtag_slave;

  //pb_cpu_to_io/m1 saved-grant jtag_uart/avalon_jtag_slave, which is an e_assign
  assign pb_cpu_to_io_m1_saved_grant_jtag_uart_avalon_jtag_slave = pb_cpu_to_io_m1_requests_jtag_uart_avalon_jtag_slave;

  //allow new arb cycle for jtag_uart/avalon_jtag_slave, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign jtag_uart_avalon_jtag_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign jtag_uart_avalon_jtag_slave_master_qreq_vector = 1;

  //jtag_uart_avalon_jtag_slave_reset_n assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_reset_n = reset_n;

  assign jtag_uart_avalon_jtag_slave_chipselect = pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave;
  //jtag_uart_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_firsttransfer = jtag_uart_avalon_jtag_slave_begins_xfer ? jtag_uart_avalon_jtag_slave_unreg_firsttransfer : jtag_uart_avalon_jtag_slave_reg_firsttransfer;

  //jtag_uart_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_unreg_firsttransfer = ~(jtag_uart_avalon_jtag_slave_slavearbiterlockenable & jtag_uart_avalon_jtag_slave_any_continuerequest);

  //jtag_uart_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_reg_firsttransfer <= 1'b1;
      else if (jtag_uart_avalon_jtag_slave_begins_xfer)
          jtag_uart_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
    end


  //jtag_uart_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_beginbursttransfer_internal = jtag_uart_avalon_jtag_slave_begins_xfer;

  //~jtag_uart_avalon_jtag_slave_read_n assignment, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_read_n = ~(pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect));

  //~jtag_uart_avalon_jtag_slave_write_n assignment, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_write_n = ~(pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect));

  assign shifted_address_to_jtag_uart_avalon_jtag_slave_from_pb_cpu_to_io_m1 = pb_cpu_to_io_m1_address_to_slave;
  //jtag_uart_avalon_jtag_slave_address mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_address = shifted_address_to_jtag_uart_avalon_jtag_slave_from_pb_cpu_to_io_m1 >> 2;

  //d1_jtag_uart_avalon_jtag_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_jtag_uart_avalon_jtag_slave_end_xfer <= 1;
      else 
        d1_jtag_uart_avalon_jtag_slave_end_xfer <= jtag_uart_avalon_jtag_slave_end_xfer;
    end


  //jtag_uart_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_waits_for_read = jtag_uart_avalon_jtag_slave_in_a_read_cycle & jtag_uart_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_in_a_read_cycle = pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = jtag_uart_avalon_jtag_slave_in_a_read_cycle;

  //jtag_uart_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_waits_for_write = jtag_uart_avalon_jtag_slave_in_a_write_cycle & jtag_uart_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_in_a_write_cycle = pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = jtag_uart_avalon_jtag_slave_in_a_write_cycle;

  assign wait_for_jtag_uart_avalon_jtag_slave_counter = 0;
  //assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //jtag_uart/avalon_jtag_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pb_cpu_to_io/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_io_m1_requests_jtag_uart_avalon_jtag_slave && (pb_cpu_to_io_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pb_cpu_to_io/m1 drove 0 on its 'burstcount' port while accessing slave jtag_uart/avalon_jtag_slave", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module led_pio_s1_arbitrator (
                               // inputs:
                                clk,
                                led_pio_s1_readdata,
                                pb_cpu_to_io_m1_address_to_slave,
                                pb_cpu_to_io_m1_burstcount,
                                pb_cpu_to_io_m1_chipselect,
                                pb_cpu_to_io_m1_latency_counter,
                                pb_cpu_to_io_m1_read,
                                pb_cpu_to_io_m1_write,
                                pb_cpu_to_io_m1_writedata,
                                reset_n,

                               // outputs:
                                d1_led_pio_s1_end_xfer,
                                led_pio_s1_address,
                                led_pio_s1_chipselect,
                                led_pio_s1_readdata_from_sa,
                                led_pio_s1_reset_n,
                                led_pio_s1_write_n,
                                led_pio_s1_writedata,
                                pb_cpu_to_io_m1_granted_led_pio_s1,
                                pb_cpu_to_io_m1_qualified_request_led_pio_s1,
                                pb_cpu_to_io_m1_read_data_valid_led_pio_s1,
                                pb_cpu_to_io_m1_requests_led_pio_s1
                             )
;

  output           d1_led_pio_s1_end_xfer;
  output  [  1: 0] led_pio_s1_address;
  output           led_pio_s1_chipselect;
  output  [ 15: 0] led_pio_s1_readdata_from_sa;
  output           led_pio_s1_reset_n;
  output           led_pio_s1_write_n;
  output  [ 15: 0] led_pio_s1_writedata;
  output           pb_cpu_to_io_m1_granted_led_pio_s1;
  output           pb_cpu_to_io_m1_qualified_request_led_pio_s1;
  output           pb_cpu_to_io_m1_read_data_valid_led_pio_s1;
  output           pb_cpu_to_io_m1_requests_led_pio_s1;
  input            clk;
  input   [ 15: 0] led_pio_s1_readdata;
  input   [ 22: 0] pb_cpu_to_io_m1_address_to_slave;
  input            pb_cpu_to_io_m1_burstcount;
  input            pb_cpu_to_io_m1_chipselect;
  input            pb_cpu_to_io_m1_latency_counter;
  input            pb_cpu_to_io_m1_read;
  input            pb_cpu_to_io_m1_write;
  input   [ 31: 0] pb_cpu_to_io_m1_writedata;
  input            reset_n;

  reg              d1_led_pio_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_led_pio_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  1: 0] led_pio_s1_address;
  wire             led_pio_s1_allgrants;
  wire             led_pio_s1_allow_new_arb_cycle;
  wire             led_pio_s1_any_bursting_master_saved_grant;
  wire             led_pio_s1_any_continuerequest;
  wire             led_pio_s1_arb_counter_enable;
  reg              led_pio_s1_arb_share_counter;
  wire             led_pio_s1_arb_share_counter_next_value;
  wire             led_pio_s1_arb_share_set_values;
  wire             led_pio_s1_beginbursttransfer_internal;
  wire             led_pio_s1_begins_xfer;
  wire             led_pio_s1_chipselect;
  wire             led_pio_s1_end_xfer;
  wire             led_pio_s1_firsttransfer;
  wire             led_pio_s1_grant_vector;
  wire             led_pio_s1_in_a_read_cycle;
  wire             led_pio_s1_in_a_write_cycle;
  wire             led_pio_s1_master_qreq_vector;
  wire             led_pio_s1_non_bursting_master_requests;
  wire    [ 15: 0] led_pio_s1_readdata_from_sa;
  reg              led_pio_s1_reg_firsttransfer;
  wire             led_pio_s1_reset_n;
  reg              led_pio_s1_slavearbiterlockenable;
  wire             led_pio_s1_slavearbiterlockenable2;
  wire             led_pio_s1_unreg_firsttransfer;
  wire             led_pio_s1_waits_for_read;
  wire             led_pio_s1_waits_for_write;
  wire             led_pio_s1_write_n;
  wire    [ 15: 0] led_pio_s1_writedata;
  wire             pb_cpu_to_io_m1_arbiterlock;
  wire             pb_cpu_to_io_m1_arbiterlock2;
  wire             pb_cpu_to_io_m1_continuerequest;
  wire             pb_cpu_to_io_m1_granted_led_pio_s1;
  wire             pb_cpu_to_io_m1_qualified_request_led_pio_s1;
  wire             pb_cpu_to_io_m1_read_data_valid_led_pio_s1;
  wire             pb_cpu_to_io_m1_requests_led_pio_s1;
  wire             pb_cpu_to_io_m1_saved_grant_led_pio_s1;
  wire    [ 22: 0] shifted_address_to_led_pio_s1_from_pb_cpu_to_io_m1;
  wire             wait_for_led_pio_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~led_pio_s1_end_xfer;
    end


  assign led_pio_s1_begins_xfer = ~d1_reasons_to_wait & ((pb_cpu_to_io_m1_qualified_request_led_pio_s1));
  //assign led_pio_s1_readdata_from_sa = led_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign led_pio_s1_readdata_from_sa = led_pio_s1_readdata;

  assign pb_cpu_to_io_m1_requests_led_pio_s1 = ({pb_cpu_to_io_m1_address_to_slave[22 : 4] , 4'b0} == 23'h4cc0) & pb_cpu_to_io_m1_chipselect;
  //led_pio_s1_arb_share_counter set values, which is an e_mux
  assign led_pio_s1_arb_share_set_values = 1;

  //led_pio_s1_non_bursting_master_requests mux, which is an e_mux
  assign led_pio_s1_non_bursting_master_requests = pb_cpu_to_io_m1_requests_led_pio_s1;

  //led_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign led_pio_s1_any_bursting_master_saved_grant = 0;

  //led_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign led_pio_s1_arb_share_counter_next_value = led_pio_s1_firsttransfer ? (led_pio_s1_arb_share_set_values - 1) : |led_pio_s1_arb_share_counter ? (led_pio_s1_arb_share_counter - 1) : 0;

  //led_pio_s1_allgrants all slave grants, which is an e_mux
  assign led_pio_s1_allgrants = |led_pio_s1_grant_vector;

  //led_pio_s1_end_xfer assignment, which is an e_assign
  assign led_pio_s1_end_xfer = ~(led_pio_s1_waits_for_read | led_pio_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_led_pio_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_led_pio_s1 = led_pio_s1_end_xfer & (~led_pio_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //led_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign led_pio_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_led_pio_s1 & led_pio_s1_allgrants) | (end_xfer_arb_share_counter_term_led_pio_s1 & ~led_pio_s1_non_bursting_master_requests);

  //led_pio_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          led_pio_s1_arb_share_counter <= 0;
      else if (led_pio_s1_arb_counter_enable)
          led_pio_s1_arb_share_counter <= led_pio_s1_arb_share_counter_next_value;
    end


  //led_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          led_pio_s1_slavearbiterlockenable <= 0;
      else if ((|led_pio_s1_master_qreq_vector & end_xfer_arb_share_counter_term_led_pio_s1) | (end_xfer_arb_share_counter_term_led_pio_s1 & ~led_pio_s1_non_bursting_master_requests))
          led_pio_s1_slavearbiterlockenable <= |led_pio_s1_arb_share_counter_next_value;
    end


  //pb_cpu_to_io/m1 led_pio/s1 arbiterlock, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock = led_pio_s1_slavearbiterlockenable & pb_cpu_to_io_m1_continuerequest;

  //led_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign led_pio_s1_slavearbiterlockenable2 = |led_pio_s1_arb_share_counter_next_value;

  //pb_cpu_to_io/m1 led_pio/s1 arbiterlock2, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock2 = led_pio_s1_slavearbiterlockenable2 & pb_cpu_to_io_m1_continuerequest;

  //led_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign led_pio_s1_any_continuerequest = 1;

  //pb_cpu_to_io_m1_continuerequest continued request, which is an e_assign
  assign pb_cpu_to_io_m1_continuerequest = 1;

  assign pb_cpu_to_io_m1_qualified_request_led_pio_s1 = pb_cpu_to_io_m1_requests_led_pio_s1 & ~(((pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ((pb_cpu_to_io_m1_latency_counter != 0))));
  //local readdatavalid pb_cpu_to_io_m1_read_data_valid_led_pio_s1, which is an e_mux
  assign pb_cpu_to_io_m1_read_data_valid_led_pio_s1 = pb_cpu_to_io_m1_granted_led_pio_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ~led_pio_s1_waits_for_read;

  //led_pio_s1_writedata mux, which is an e_mux
  assign led_pio_s1_writedata = pb_cpu_to_io_m1_writedata;

  //master is always granted when requested
  assign pb_cpu_to_io_m1_granted_led_pio_s1 = pb_cpu_to_io_m1_qualified_request_led_pio_s1;

  //pb_cpu_to_io/m1 saved-grant led_pio/s1, which is an e_assign
  assign pb_cpu_to_io_m1_saved_grant_led_pio_s1 = pb_cpu_to_io_m1_requests_led_pio_s1;

  //allow new arb cycle for led_pio/s1, which is an e_assign
  assign led_pio_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign led_pio_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign led_pio_s1_master_qreq_vector = 1;

  //led_pio_s1_reset_n assignment, which is an e_assign
  assign led_pio_s1_reset_n = reset_n;

  assign led_pio_s1_chipselect = pb_cpu_to_io_m1_granted_led_pio_s1;
  //led_pio_s1_firsttransfer first transaction, which is an e_assign
  assign led_pio_s1_firsttransfer = led_pio_s1_begins_xfer ? led_pio_s1_unreg_firsttransfer : led_pio_s1_reg_firsttransfer;

  //led_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign led_pio_s1_unreg_firsttransfer = ~(led_pio_s1_slavearbiterlockenable & led_pio_s1_any_continuerequest);

  //led_pio_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          led_pio_s1_reg_firsttransfer <= 1'b1;
      else if (led_pio_s1_begins_xfer)
          led_pio_s1_reg_firsttransfer <= led_pio_s1_unreg_firsttransfer;
    end


  //led_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign led_pio_s1_beginbursttransfer_internal = led_pio_s1_begins_xfer;

  //~led_pio_s1_write_n assignment, which is an e_mux
  assign led_pio_s1_write_n = ~(pb_cpu_to_io_m1_granted_led_pio_s1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect));

  assign shifted_address_to_led_pio_s1_from_pb_cpu_to_io_m1 = pb_cpu_to_io_m1_address_to_slave;
  //led_pio_s1_address mux, which is an e_mux
  assign led_pio_s1_address = shifted_address_to_led_pio_s1_from_pb_cpu_to_io_m1 >> 2;

  //d1_led_pio_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_led_pio_s1_end_xfer <= 1;
      else 
        d1_led_pio_s1_end_xfer <= led_pio_s1_end_xfer;
    end


  //led_pio_s1_waits_for_read in a cycle, which is an e_mux
  assign led_pio_s1_waits_for_read = led_pio_s1_in_a_read_cycle & led_pio_s1_begins_xfer;

  //led_pio_s1_in_a_read_cycle assignment, which is an e_assign
  assign led_pio_s1_in_a_read_cycle = pb_cpu_to_io_m1_granted_led_pio_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = led_pio_s1_in_a_read_cycle;

  //led_pio_s1_waits_for_write in a cycle, which is an e_mux
  assign led_pio_s1_waits_for_write = led_pio_s1_in_a_write_cycle & 0;

  //led_pio_s1_in_a_write_cycle assignment, which is an e_assign
  assign led_pio_s1_in_a_write_cycle = pb_cpu_to_io_m1_granted_led_pio_s1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = led_pio_s1_in_a_write_cycle;

  assign wait_for_led_pio_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //led_pio/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pb_cpu_to_io/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_io_m1_requests_led_pio_s1 && (pb_cpu_to_io_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pb_cpu_to_io/m1 drove 0 on its 'burstcount' port while accessing slave led_pio/s1", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_pb_cpu_to_ddr3_top_s1_module (
                                                                      // inputs:
                                                                       clear_fifo,
                                                                       clk,
                                                                       data_in,
                                                                       read,
                                                                       reset_n,
                                                                       sync_reset,
                                                                       write,

                                                                      // outputs:
                                                                       data_out,
                                                                       empty,
                                                                       fifo_contains_ones_n,
                                                                       full
                                                                    )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  wire             full_34;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_33;
  assign empty = !full_0;
  assign full_34 = 0;
  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    0;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_instruction_master_to_pb_cpu_to_ddr3_top_s1_module (
                                                                             // inputs:
                                                                              clear_fifo,
                                                                              clk,
                                                                              data_in,
                                                                              read,
                                                                              reset_n,
                                                                              sync_reset,
                                                                              write,

                                                                             // outputs:
                                                                              data_out,
                                                                              empty,
                                                                              fifo_contains_ones_n,
                                                                              full
                                                                           )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  wire             full_34;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_33;
  assign empty = !full_0;
  assign full_34 = 0;
  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    0;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pb_cpu_to_ddr3_top_s1_arbitrator (
                                          // inputs:
                                           clk,
                                           cpu_data_master_address_to_slave,
                                           cpu_data_master_byteenable,
                                           cpu_data_master_debugaccess,
                                           cpu_data_master_latency_counter,
                                           cpu_data_master_read,
                                           cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register,
                                           cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register,
                                           cpu_data_master_write,
                                           cpu_data_master_writedata,
                                           cpu_instruction_master_address_to_slave,
                                           cpu_instruction_master_latency_counter,
                                           cpu_instruction_master_read,
                                           cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register,
                                           pb_cpu_to_ddr3_top_s1_endofpacket,
                                           pb_cpu_to_ddr3_top_s1_readdata,
                                           pb_cpu_to_ddr3_top_s1_readdatavalid,
                                           pb_cpu_to_ddr3_top_s1_waitrequest,
                                           reset_n,

                                          // outputs:
                                           cpu_data_master_granted_pb_cpu_to_ddr3_top_s1,
                                           cpu_data_master_qualified_request_pb_cpu_to_ddr3_top_s1,
                                           cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1,
                                           cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register,
                                           cpu_data_master_requests_pb_cpu_to_ddr3_top_s1,
                                           cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1,
                                           cpu_instruction_master_qualified_request_pb_cpu_to_ddr3_top_s1,
                                           cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1,
                                           cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register,
                                           cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1,
                                           d1_pb_cpu_to_ddr3_top_s1_end_xfer,
                                           pb_cpu_to_ddr3_top_s1_address,
                                           pb_cpu_to_ddr3_top_s1_arbiterlock,
                                           pb_cpu_to_ddr3_top_s1_arbiterlock2,
                                           pb_cpu_to_ddr3_top_s1_burstcount,
                                           pb_cpu_to_ddr3_top_s1_byteenable,
                                           pb_cpu_to_ddr3_top_s1_chipselect,
                                           pb_cpu_to_ddr3_top_s1_debugaccess,
                                           pb_cpu_to_ddr3_top_s1_endofpacket_from_sa,
                                           pb_cpu_to_ddr3_top_s1_nativeaddress,
                                           pb_cpu_to_ddr3_top_s1_read,
                                           pb_cpu_to_ddr3_top_s1_readdata_from_sa,
                                           pb_cpu_to_ddr3_top_s1_reset_n,
                                           pb_cpu_to_ddr3_top_s1_waitrequest_from_sa,
                                           pb_cpu_to_ddr3_top_s1_write,
                                           pb_cpu_to_ddr3_top_s1_writedata
                                        )
;

  output           cpu_data_master_granted_pb_cpu_to_ddr3_top_s1;
  output           cpu_data_master_qualified_request_pb_cpu_to_ddr3_top_s1;
  output           cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1;
  output           cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register;
  output           cpu_data_master_requests_pb_cpu_to_ddr3_top_s1;
  output           cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1;
  output           cpu_instruction_master_qualified_request_pb_cpu_to_ddr3_top_s1;
  output           cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1;
  output           cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register;
  output           cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1;
  output           d1_pb_cpu_to_ddr3_top_s1_end_xfer;
  output  [ 24: 0] pb_cpu_to_ddr3_top_s1_address;
  output           pb_cpu_to_ddr3_top_s1_arbiterlock;
  output           pb_cpu_to_ddr3_top_s1_arbiterlock2;
  output           pb_cpu_to_ddr3_top_s1_burstcount;
  output  [  3: 0] pb_cpu_to_ddr3_top_s1_byteenable;
  output           pb_cpu_to_ddr3_top_s1_chipselect;
  output           pb_cpu_to_ddr3_top_s1_debugaccess;
  output           pb_cpu_to_ddr3_top_s1_endofpacket_from_sa;
  output  [ 24: 0] pb_cpu_to_ddr3_top_s1_nativeaddress;
  output           pb_cpu_to_ddr3_top_s1_read;
  output  [ 31: 0] pb_cpu_to_ddr3_top_s1_readdata_from_sa;
  output           pb_cpu_to_ddr3_top_s1_reset_n;
  output           pb_cpu_to_ddr3_top_s1_waitrequest_from_sa;
  output           pb_cpu_to_ddr3_top_s1_write;
  output  [ 31: 0] pb_cpu_to_ddr3_top_s1_writedata;
  input            clk;
  input   [ 28: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register;
  input            cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 28: 0] cpu_instruction_master_address_to_slave;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register;
  input            pb_cpu_to_ddr3_top_s1_endofpacket;
  input   [ 31: 0] pb_cpu_to_ddr3_top_s1_readdata;
  input            pb_cpu_to_ddr3_top_s1_readdatavalid;
  input            pb_cpu_to_ddr3_top_s1_waitrequest;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_pb_cpu_to_ddr3_top_s1;
  wire             cpu_data_master_qualified_request_pb_cpu_to_ddr3_top_s1;
  wire             cpu_data_master_rdv_fifo_empty_pb_cpu_to_ddr3_top_s1;
  wire             cpu_data_master_rdv_fifo_output_from_pb_cpu_to_ddr3_top_s1;
  wire             cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1;
  wire             cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register;
  wire             cpu_data_master_requests_pb_cpu_to_ddr3_top_s1;
  wire             cpu_data_master_saved_grant_pb_cpu_to_ddr3_top_s1;
  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1;
  wire             cpu_instruction_master_qualified_request_pb_cpu_to_ddr3_top_s1;
  wire             cpu_instruction_master_rdv_fifo_empty_pb_cpu_to_ddr3_top_s1;
  wire             cpu_instruction_master_rdv_fifo_output_from_pb_cpu_to_ddr3_top_s1;
  wire             cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1;
  wire             cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register;
  wire             cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1;
  wire             cpu_instruction_master_saved_grant_pb_cpu_to_ddr3_top_s1;
  reg              d1_pb_cpu_to_ddr3_top_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_pb_cpu_to_ddr3_top_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_data_master_granted_slave_pb_cpu_to_ddr3_top_s1;
  reg              last_cycle_cpu_instruction_master_granted_slave_pb_cpu_to_ddr3_top_s1;
  wire    [ 24: 0] pb_cpu_to_ddr3_top_s1_address;
  wire             pb_cpu_to_ddr3_top_s1_allgrants;
  wire             pb_cpu_to_ddr3_top_s1_allow_new_arb_cycle;
  wire             pb_cpu_to_ddr3_top_s1_any_bursting_master_saved_grant;
  wire             pb_cpu_to_ddr3_top_s1_any_continuerequest;
  reg     [  1: 0] pb_cpu_to_ddr3_top_s1_arb_addend;
  wire             pb_cpu_to_ddr3_top_s1_arb_counter_enable;
  reg     [  3: 0] pb_cpu_to_ddr3_top_s1_arb_share_counter;
  wire    [  3: 0] pb_cpu_to_ddr3_top_s1_arb_share_counter_next_value;
  wire    [  3: 0] pb_cpu_to_ddr3_top_s1_arb_share_set_values;
  wire    [  1: 0] pb_cpu_to_ddr3_top_s1_arb_winner;
  wire             pb_cpu_to_ddr3_top_s1_arbiterlock;
  wire             pb_cpu_to_ddr3_top_s1_arbiterlock2;
  wire             pb_cpu_to_ddr3_top_s1_arbitration_holdoff_internal;
  wire             pb_cpu_to_ddr3_top_s1_beginbursttransfer_internal;
  wire             pb_cpu_to_ddr3_top_s1_begins_xfer;
  wire             pb_cpu_to_ddr3_top_s1_burstcount;
  wire    [  3: 0] pb_cpu_to_ddr3_top_s1_byteenable;
  wire             pb_cpu_to_ddr3_top_s1_chipselect;
  wire    [  3: 0] pb_cpu_to_ddr3_top_s1_chosen_master_double_vector;
  wire    [  1: 0] pb_cpu_to_ddr3_top_s1_chosen_master_rot_left;
  wire             pb_cpu_to_ddr3_top_s1_debugaccess;
  wire             pb_cpu_to_ddr3_top_s1_end_xfer;
  wire             pb_cpu_to_ddr3_top_s1_endofpacket_from_sa;
  wire             pb_cpu_to_ddr3_top_s1_firsttransfer;
  wire    [  1: 0] pb_cpu_to_ddr3_top_s1_grant_vector;
  wire             pb_cpu_to_ddr3_top_s1_in_a_read_cycle;
  wire             pb_cpu_to_ddr3_top_s1_in_a_write_cycle;
  wire    [  1: 0] pb_cpu_to_ddr3_top_s1_master_qreq_vector;
  wire             pb_cpu_to_ddr3_top_s1_move_on_to_next_transaction;
  wire    [ 24: 0] pb_cpu_to_ddr3_top_s1_nativeaddress;
  wire             pb_cpu_to_ddr3_top_s1_non_bursting_master_requests;
  wire             pb_cpu_to_ddr3_top_s1_read;
  wire    [ 31: 0] pb_cpu_to_ddr3_top_s1_readdata_from_sa;
  wire             pb_cpu_to_ddr3_top_s1_readdatavalid_from_sa;
  reg              pb_cpu_to_ddr3_top_s1_reg_firsttransfer;
  wire             pb_cpu_to_ddr3_top_s1_reset_n;
  reg     [  1: 0] pb_cpu_to_ddr3_top_s1_saved_chosen_master_vector;
  reg              pb_cpu_to_ddr3_top_s1_slavearbiterlockenable;
  wire             pb_cpu_to_ddr3_top_s1_slavearbiterlockenable2;
  wire             pb_cpu_to_ddr3_top_s1_unreg_firsttransfer;
  wire             pb_cpu_to_ddr3_top_s1_waitrequest_from_sa;
  wire             pb_cpu_to_ddr3_top_s1_waits_for_read;
  wire             pb_cpu_to_ddr3_top_s1_waits_for_write;
  wire             pb_cpu_to_ddr3_top_s1_write;
  wire    [ 31: 0] pb_cpu_to_ddr3_top_s1_writedata;
  wire    [ 28: 0] shifted_address_to_pb_cpu_to_ddr3_top_s1_from_cpu_data_master;
  wire    [ 28: 0] shifted_address_to_pb_cpu_to_ddr3_top_s1_from_cpu_instruction_master;
  wire             wait_for_pb_cpu_to_ddr3_top_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~pb_cpu_to_ddr3_top_s1_end_xfer;
    end


  assign pb_cpu_to_ddr3_top_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_pb_cpu_to_ddr3_top_s1 | cpu_instruction_master_qualified_request_pb_cpu_to_ddr3_top_s1));
  //assign pb_cpu_to_ddr3_top_s1_readdatavalid_from_sa = pb_cpu_to_ddr3_top_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_readdatavalid_from_sa = pb_cpu_to_ddr3_top_s1_readdatavalid;

  //assign pb_cpu_to_ddr3_top_s1_readdata_from_sa = pb_cpu_to_ddr3_top_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_readdata_from_sa = pb_cpu_to_ddr3_top_s1_readdata;

  assign cpu_data_master_requests_pb_cpu_to_ddr3_top_s1 = ({cpu_data_master_address_to_slave[28 : 27] , 27'b0} == 29'h10000000) & (cpu_data_master_read | cpu_data_master_write);
  //assign pb_cpu_to_ddr3_top_s1_waitrequest_from_sa = pb_cpu_to_ddr3_top_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_waitrequest_from_sa = pb_cpu_to_ddr3_top_s1_waitrequest;

  //pb_cpu_to_ddr3_top_s1_arb_share_counter set values, which is an e_mux
  assign pb_cpu_to_ddr3_top_s1_arb_share_set_values = (cpu_data_master_granted_pb_cpu_to_ddr3_top_s1)? 8 :
    (cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1)? 8 :
    (cpu_data_master_granted_pb_cpu_to_ddr3_top_s1)? 8 :
    (cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1)? 8 :
    (cpu_data_master_granted_pb_cpu_to_ddr3_top_s1)? 8 :
    (cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1)? 8 :
    1;

  //pb_cpu_to_ddr3_top_s1_non_bursting_master_requests mux, which is an e_mux
  assign pb_cpu_to_ddr3_top_s1_non_bursting_master_requests = cpu_data_master_requests_pb_cpu_to_ddr3_top_s1 |
    cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1 |
    cpu_data_master_requests_pb_cpu_to_ddr3_top_s1 |
    cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1 |
    cpu_data_master_requests_pb_cpu_to_ddr3_top_s1 |
    cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1;

  //pb_cpu_to_ddr3_top_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign pb_cpu_to_ddr3_top_s1_any_bursting_master_saved_grant = 0;

  //pb_cpu_to_ddr3_top_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_arb_share_counter_next_value = pb_cpu_to_ddr3_top_s1_firsttransfer ? (pb_cpu_to_ddr3_top_s1_arb_share_set_values - 1) : |pb_cpu_to_ddr3_top_s1_arb_share_counter ? (pb_cpu_to_ddr3_top_s1_arb_share_counter - 1) : 0;

  //pb_cpu_to_ddr3_top_s1_allgrants all slave grants, which is an e_mux
  assign pb_cpu_to_ddr3_top_s1_allgrants = (|pb_cpu_to_ddr3_top_s1_grant_vector) |
    (|pb_cpu_to_ddr3_top_s1_grant_vector) |
    (|pb_cpu_to_ddr3_top_s1_grant_vector) |
    (|pb_cpu_to_ddr3_top_s1_grant_vector) |
    (|pb_cpu_to_ddr3_top_s1_grant_vector) |
    (|pb_cpu_to_ddr3_top_s1_grant_vector);

  //pb_cpu_to_ddr3_top_s1_end_xfer assignment, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_end_xfer = ~(pb_cpu_to_ddr3_top_s1_waits_for_read | pb_cpu_to_ddr3_top_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_pb_cpu_to_ddr3_top_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_pb_cpu_to_ddr3_top_s1 = pb_cpu_to_ddr3_top_s1_end_xfer & (~pb_cpu_to_ddr3_top_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //pb_cpu_to_ddr3_top_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_pb_cpu_to_ddr3_top_s1 & pb_cpu_to_ddr3_top_s1_allgrants) | (end_xfer_arb_share_counter_term_pb_cpu_to_ddr3_top_s1 & ~pb_cpu_to_ddr3_top_s1_non_bursting_master_requests);

  //pb_cpu_to_ddr3_top_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_ddr3_top_s1_arb_share_counter <= 0;
      else if (pb_cpu_to_ddr3_top_s1_arb_counter_enable)
          pb_cpu_to_ddr3_top_s1_arb_share_counter <= pb_cpu_to_ddr3_top_s1_arb_share_counter_next_value;
    end


  //pb_cpu_to_ddr3_top_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_ddr3_top_s1_slavearbiterlockenable <= 0;
      else if ((|pb_cpu_to_ddr3_top_s1_master_qreq_vector & end_xfer_arb_share_counter_term_pb_cpu_to_ddr3_top_s1) | (end_xfer_arb_share_counter_term_pb_cpu_to_ddr3_top_s1 & ~pb_cpu_to_ddr3_top_s1_non_bursting_master_requests))
          pb_cpu_to_ddr3_top_s1_slavearbiterlockenable <= |pb_cpu_to_ddr3_top_s1_arb_share_counter_next_value;
    end


  //cpu/data_master pb_cpu_to_ddr3_top/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = pb_cpu_to_ddr3_top_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //pb_cpu_to_ddr3_top_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_slavearbiterlockenable2 = |pb_cpu_to_ddr3_top_s1_arb_share_counter_next_value;

  //cpu/data_master pb_cpu_to_ddr3_top/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = pb_cpu_to_ddr3_top_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //cpu/instruction_master pb_cpu_to_ddr3_top/s1 arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = pb_cpu_to_ddr3_top_s1_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //cpu/instruction_master pb_cpu_to_ddr3_top/s1 arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = pb_cpu_to_ddr3_top_s1_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //cpu/instruction_master granted pb_cpu_to_ddr3_top/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_instruction_master_granted_slave_pb_cpu_to_ddr3_top_s1 <= 0;
      else 
        last_cycle_cpu_instruction_master_granted_slave_pb_cpu_to_ddr3_top_s1 <= cpu_instruction_master_saved_grant_pb_cpu_to_ddr3_top_s1 ? 1 : (pb_cpu_to_ddr3_top_s1_arbitration_holdoff_internal | ~cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1) ? 0 : last_cycle_cpu_instruction_master_granted_slave_pb_cpu_to_ddr3_top_s1;
    end


  //cpu_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_instruction_master_continuerequest = last_cycle_cpu_instruction_master_granted_slave_pb_cpu_to_ddr3_top_s1 & cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1;

  //pb_cpu_to_ddr3_top_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign pb_cpu_to_ddr3_top_s1_any_continuerequest = cpu_instruction_master_continuerequest |
    cpu_data_master_continuerequest;

  assign cpu_data_master_qualified_request_pb_cpu_to_ddr3_top_s1 = cpu_data_master_requests_pb_cpu_to_ddr3_top_s1 & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register) | (|cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register))) | cpu_instruction_master_arbiterlock);
  //unique name for pb_cpu_to_ddr3_top_s1_move_on_to_next_transaction, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_move_on_to_next_transaction = pb_cpu_to_ddr3_top_s1_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_pb_cpu_to_ddr3_top_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_pb_cpu_to_ddr3_top_s1_module rdv_fifo_for_cpu_data_master_to_pb_cpu_to_ddr3_top_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_pb_cpu_to_ddr3_top_s1),
      .data_out             (cpu_data_master_rdv_fifo_output_from_pb_cpu_to_ddr3_top_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_pb_cpu_to_ddr3_top_s1),
      .full                 (),
      .read                 (pb_cpu_to_ddr3_top_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~pb_cpu_to_ddr3_top_s1_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register = ~cpu_data_master_rdv_fifo_empty_pb_cpu_to_ddr3_top_s1;
  //local readdatavalid cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1 = (pb_cpu_to_ddr3_top_s1_readdatavalid_from_sa & cpu_data_master_rdv_fifo_output_from_pb_cpu_to_ddr3_top_s1) & ~ cpu_data_master_rdv_fifo_empty_pb_cpu_to_ddr3_top_s1;

  //pb_cpu_to_ddr3_top_s1_writedata mux, which is an e_mux
  assign pb_cpu_to_ddr3_top_s1_writedata = cpu_data_master_writedata;

  //assign pb_cpu_to_ddr3_top_s1_endofpacket_from_sa = pb_cpu_to_ddr3_top_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_endofpacket_from_sa = pb_cpu_to_ddr3_top_s1_endofpacket;

  assign cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1 = (({cpu_instruction_master_address_to_slave[28 : 27] , 27'b0} == 29'h10000000) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //cpu/data_master granted pb_cpu_to_ddr3_top/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_data_master_granted_slave_pb_cpu_to_ddr3_top_s1 <= 0;
      else 
        last_cycle_cpu_data_master_granted_slave_pb_cpu_to_ddr3_top_s1 <= cpu_data_master_saved_grant_pb_cpu_to_ddr3_top_s1 ? 1 : (pb_cpu_to_ddr3_top_s1_arbitration_holdoff_internal | ~cpu_data_master_requests_pb_cpu_to_ddr3_top_s1) ? 0 : last_cycle_cpu_data_master_granted_slave_pb_cpu_to_ddr3_top_s1;
    end


  //cpu_data_master_continuerequest continued request, which is an e_mux
  assign cpu_data_master_continuerequest = last_cycle_cpu_data_master_granted_slave_pb_cpu_to_ddr3_top_s1 & cpu_data_master_requests_pb_cpu_to_ddr3_top_s1;

  assign cpu_instruction_master_qualified_request_pb_cpu_to_ddr3_top_s1 = cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1 & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (1 < cpu_instruction_master_latency_counter) | (|cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register))) | cpu_data_master_arbiterlock);
  //rdv_fifo_for_cpu_instruction_master_to_pb_cpu_to_ddr3_top_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_pb_cpu_to_ddr3_top_s1_module rdv_fifo_for_cpu_instruction_master_to_pb_cpu_to_ddr3_top_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1),
      .data_out             (cpu_instruction_master_rdv_fifo_output_from_pb_cpu_to_ddr3_top_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_instruction_master_rdv_fifo_empty_pb_cpu_to_ddr3_top_s1),
      .full                 (),
      .read                 (pb_cpu_to_ddr3_top_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~pb_cpu_to_ddr3_top_s1_waits_for_read)
    );

  assign cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register = ~cpu_instruction_master_rdv_fifo_empty_pb_cpu_to_ddr3_top_s1;
  //local readdatavalid cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1, which is an e_mux
  assign cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1 = (pb_cpu_to_ddr3_top_s1_readdatavalid_from_sa & cpu_instruction_master_rdv_fifo_output_from_pb_cpu_to_ddr3_top_s1) & ~ cpu_instruction_master_rdv_fifo_empty_pb_cpu_to_ddr3_top_s1;

  //allow new arb cycle for pb_cpu_to_ddr3_top/s1, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_allow_new_arb_cycle = ~cpu_data_master_arbiterlock & ~cpu_instruction_master_arbiterlock;

  //cpu/instruction_master assignment into master qualified-requests vector for pb_cpu_to_ddr3_top/s1, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_master_qreq_vector[0] = cpu_instruction_master_qualified_request_pb_cpu_to_ddr3_top_s1;

  //cpu/instruction_master grant pb_cpu_to_ddr3_top/s1, which is an e_assign
  assign cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1 = pb_cpu_to_ddr3_top_s1_grant_vector[0];

  //cpu/instruction_master saved-grant pb_cpu_to_ddr3_top/s1, which is an e_assign
  assign cpu_instruction_master_saved_grant_pb_cpu_to_ddr3_top_s1 = pb_cpu_to_ddr3_top_s1_arb_winner[0] && cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1;

  //cpu/data_master assignment into master qualified-requests vector for pb_cpu_to_ddr3_top/s1, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_master_qreq_vector[1] = cpu_data_master_qualified_request_pb_cpu_to_ddr3_top_s1;

  //cpu/data_master grant pb_cpu_to_ddr3_top/s1, which is an e_assign
  assign cpu_data_master_granted_pb_cpu_to_ddr3_top_s1 = pb_cpu_to_ddr3_top_s1_grant_vector[1];

  //cpu/data_master saved-grant pb_cpu_to_ddr3_top/s1, which is an e_assign
  assign cpu_data_master_saved_grant_pb_cpu_to_ddr3_top_s1 = pb_cpu_to_ddr3_top_s1_arb_winner[1] && cpu_data_master_requests_pb_cpu_to_ddr3_top_s1;

  //pb_cpu_to_ddr3_top/s1 chosen-master double-vector, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_chosen_master_double_vector = {pb_cpu_to_ddr3_top_s1_master_qreq_vector, pb_cpu_to_ddr3_top_s1_master_qreq_vector} & ({~pb_cpu_to_ddr3_top_s1_master_qreq_vector, ~pb_cpu_to_ddr3_top_s1_master_qreq_vector} + pb_cpu_to_ddr3_top_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign pb_cpu_to_ddr3_top_s1_arb_winner = (pb_cpu_to_ddr3_top_s1_allow_new_arb_cycle & | pb_cpu_to_ddr3_top_s1_grant_vector) ? pb_cpu_to_ddr3_top_s1_grant_vector : pb_cpu_to_ddr3_top_s1_saved_chosen_master_vector;

  //saved pb_cpu_to_ddr3_top_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_ddr3_top_s1_saved_chosen_master_vector <= 0;
      else if (pb_cpu_to_ddr3_top_s1_allow_new_arb_cycle)
          pb_cpu_to_ddr3_top_s1_saved_chosen_master_vector <= |pb_cpu_to_ddr3_top_s1_grant_vector ? pb_cpu_to_ddr3_top_s1_grant_vector : pb_cpu_to_ddr3_top_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign pb_cpu_to_ddr3_top_s1_grant_vector = {(pb_cpu_to_ddr3_top_s1_chosen_master_double_vector[1] | pb_cpu_to_ddr3_top_s1_chosen_master_double_vector[3]),
    (pb_cpu_to_ddr3_top_s1_chosen_master_double_vector[0] | pb_cpu_to_ddr3_top_s1_chosen_master_double_vector[2])};

  //pb_cpu_to_ddr3_top/s1 chosen master rotated left, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_chosen_master_rot_left = (pb_cpu_to_ddr3_top_s1_arb_winner << 1) ? (pb_cpu_to_ddr3_top_s1_arb_winner << 1) : 1;

  //pb_cpu_to_ddr3_top/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_ddr3_top_s1_arb_addend <= 1;
      else if (|pb_cpu_to_ddr3_top_s1_grant_vector)
          pb_cpu_to_ddr3_top_s1_arb_addend <= pb_cpu_to_ddr3_top_s1_end_xfer? pb_cpu_to_ddr3_top_s1_chosen_master_rot_left : pb_cpu_to_ddr3_top_s1_grant_vector;
    end


  //pb_cpu_to_ddr3_top_s1_reset_n assignment, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_reset_n = reset_n;

  assign pb_cpu_to_ddr3_top_s1_chipselect = cpu_data_master_granted_pb_cpu_to_ddr3_top_s1 | cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1;
  //pb_cpu_to_ddr3_top_s1_firsttransfer first transaction, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_firsttransfer = pb_cpu_to_ddr3_top_s1_begins_xfer ? pb_cpu_to_ddr3_top_s1_unreg_firsttransfer : pb_cpu_to_ddr3_top_s1_reg_firsttransfer;

  //pb_cpu_to_ddr3_top_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_unreg_firsttransfer = ~(pb_cpu_to_ddr3_top_s1_slavearbiterlockenable & pb_cpu_to_ddr3_top_s1_any_continuerequest);

  //pb_cpu_to_ddr3_top_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_ddr3_top_s1_reg_firsttransfer <= 1'b1;
      else if (pb_cpu_to_ddr3_top_s1_begins_xfer)
          pb_cpu_to_ddr3_top_s1_reg_firsttransfer <= pb_cpu_to_ddr3_top_s1_unreg_firsttransfer;
    end


  //pb_cpu_to_ddr3_top_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_beginbursttransfer_internal = pb_cpu_to_ddr3_top_s1_begins_xfer;

  //pb_cpu_to_ddr3_top_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_arbitration_holdoff_internal = pb_cpu_to_ddr3_top_s1_begins_xfer & pb_cpu_to_ddr3_top_s1_firsttransfer;

  //pb_cpu_to_ddr3_top_s1_read assignment, which is an e_mux
  assign pb_cpu_to_ddr3_top_s1_read = (cpu_data_master_granted_pb_cpu_to_ddr3_top_s1 & cpu_data_master_read) | (cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1 & cpu_instruction_master_read);

  //pb_cpu_to_ddr3_top_s1_write assignment, which is an e_mux
  assign pb_cpu_to_ddr3_top_s1_write = cpu_data_master_granted_pb_cpu_to_ddr3_top_s1 & cpu_data_master_write;

  assign shifted_address_to_pb_cpu_to_ddr3_top_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //pb_cpu_to_ddr3_top_s1_address mux, which is an e_mux
  assign pb_cpu_to_ddr3_top_s1_address = (cpu_data_master_granted_pb_cpu_to_ddr3_top_s1)? (shifted_address_to_pb_cpu_to_ddr3_top_s1_from_cpu_data_master >> 2) :
    (shifted_address_to_pb_cpu_to_ddr3_top_s1_from_cpu_instruction_master >> 2);

  assign shifted_address_to_pb_cpu_to_ddr3_top_s1_from_cpu_instruction_master = cpu_instruction_master_address_to_slave;
  //slaveid pb_cpu_to_ddr3_top_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign pb_cpu_to_ddr3_top_s1_nativeaddress = (cpu_data_master_granted_pb_cpu_to_ddr3_top_s1)? (cpu_data_master_address_to_slave >> 2) :
    (cpu_instruction_master_address_to_slave >> 2);

  //d1_pb_cpu_to_ddr3_top_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_pb_cpu_to_ddr3_top_s1_end_xfer <= 1;
      else 
        d1_pb_cpu_to_ddr3_top_s1_end_xfer <= pb_cpu_to_ddr3_top_s1_end_xfer;
    end


  //pb_cpu_to_ddr3_top_s1_waits_for_read in a cycle, which is an e_mux
  assign pb_cpu_to_ddr3_top_s1_waits_for_read = pb_cpu_to_ddr3_top_s1_in_a_read_cycle & pb_cpu_to_ddr3_top_s1_waitrequest_from_sa;

  //pb_cpu_to_ddr3_top_s1_in_a_read_cycle assignment, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_in_a_read_cycle = (cpu_data_master_granted_pb_cpu_to_ddr3_top_s1 & cpu_data_master_read) | (cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1 & cpu_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = pb_cpu_to_ddr3_top_s1_in_a_read_cycle;

  //pb_cpu_to_ddr3_top_s1_waits_for_write in a cycle, which is an e_mux
  assign pb_cpu_to_ddr3_top_s1_waits_for_write = pb_cpu_to_ddr3_top_s1_in_a_write_cycle & pb_cpu_to_ddr3_top_s1_waitrequest_from_sa;

  //pb_cpu_to_ddr3_top_s1_in_a_write_cycle assignment, which is an e_assign
  assign pb_cpu_to_ddr3_top_s1_in_a_write_cycle = cpu_data_master_granted_pb_cpu_to_ddr3_top_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = pb_cpu_to_ddr3_top_s1_in_a_write_cycle;

  assign wait_for_pb_cpu_to_ddr3_top_s1_counter = 0;
  //pb_cpu_to_ddr3_top_s1_byteenable byte enable port mux, which is an e_mux
  assign pb_cpu_to_ddr3_top_s1_byteenable = (cpu_data_master_granted_pb_cpu_to_ddr3_top_s1)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign pb_cpu_to_ddr3_top_s1_burstcount = 1;

  //pb_cpu_to_ddr3_top/s1 arbiterlock assigned from _handle_arbiterlock, which is an e_mux
  assign pb_cpu_to_ddr3_top_s1_arbiterlock = (cpu_data_master_arbiterlock)? cpu_data_master_arbiterlock :
    cpu_instruction_master_arbiterlock;

  //pb_cpu_to_ddr3_top/s1 arbiterlock2 assigned from _handle_arbiterlock2, which is an e_mux
  assign pb_cpu_to_ddr3_top_s1_arbiterlock2 = (cpu_data_master_arbiterlock2)? cpu_data_master_arbiterlock2 :
    cpu_instruction_master_arbiterlock2;

  //debugaccess mux, which is an e_mux
  assign pb_cpu_to_ddr3_top_s1_debugaccess = (cpu_data_master_granted_pb_cpu_to_ddr3_top_s1)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pb_cpu_to_ddr3_top/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_granted_pb_cpu_to_ddr3_top_s1 + cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_saved_grant_pb_cpu_to_ddr3_top_s1 + cpu_instruction_master_saved_grant_pb_cpu_to_ddr3_top_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo_module (
                                                                      // inputs:
                                                                       clear_fifo,
                                                                       clk,
                                                                       data_in,
                                                                       read,
                                                                       reset_n,
                                                                       sync_reset,
                                                                       write,

                                                                      // outputs:
                                                                       data_out,
                                                                       empty,
                                                                       fifo_contains_ones_n,
                                                                       full
                                                                    )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  wire             full_32;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_31;
  assign empty = !full_0;
  assign full_32 = 0;
  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    0;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pb_cpu_to_ddr3_top_m1_arbitrator (
                                          // inputs:
                                           clk,
                                           d1_ddr3_top_s1_end_xfer,
                                           ddr3_top_s1_readdata_from_sa,
                                           ddr3_top_s1_waitrequest_n_from_sa,
                                           pb_cpu_to_ddr3_top_m1_address,
                                           pb_cpu_to_ddr3_top_m1_burstcount,
                                           pb_cpu_to_ddr3_top_m1_byteenable,
                                           pb_cpu_to_ddr3_top_m1_chipselect,
                                           pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1,
                                           pb_cpu_to_ddr3_top_m1_qualified_request_ddr3_top_s1,
                                           pb_cpu_to_ddr3_top_m1_read,
                                           pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1,
                                           pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register,
                                           pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1,
                                           pb_cpu_to_ddr3_top_m1_write,
                                           pb_cpu_to_ddr3_top_m1_writedata,
                                           reset_n,

                                          // outputs:
                                           pb_cpu_to_ddr3_top_m1_address_to_slave,
                                           pb_cpu_to_ddr3_top_m1_latency_counter,
                                           pb_cpu_to_ddr3_top_m1_readdata,
                                           pb_cpu_to_ddr3_top_m1_readdatavalid,
                                           pb_cpu_to_ddr3_top_m1_waitrequest
                                        )
;

  output  [ 26: 0] pb_cpu_to_ddr3_top_m1_address_to_slave;
  output           pb_cpu_to_ddr3_top_m1_latency_counter;
  output  [ 31: 0] pb_cpu_to_ddr3_top_m1_readdata;
  output           pb_cpu_to_ddr3_top_m1_readdatavalid;
  output           pb_cpu_to_ddr3_top_m1_waitrequest;
  input            clk;
  input            d1_ddr3_top_s1_end_xfer;
  input   [ 63: 0] ddr3_top_s1_readdata_from_sa;
  input            ddr3_top_s1_waitrequest_n_from_sa;
  input   [ 26: 0] pb_cpu_to_ddr3_top_m1_address;
  input            pb_cpu_to_ddr3_top_m1_burstcount;
  input   [  3: 0] pb_cpu_to_ddr3_top_m1_byteenable;
  input            pb_cpu_to_ddr3_top_m1_chipselect;
  input            pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1;
  input            pb_cpu_to_ddr3_top_m1_qualified_request_ddr3_top_s1;
  input            pb_cpu_to_ddr3_top_m1_read;
  input            pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1;
  input            pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register;
  input            pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1;
  input            pb_cpu_to_ddr3_top_m1_write;
  input   [ 31: 0] pb_cpu_to_ddr3_top_m1_writedata;
  input            reset_n;

  reg              active_and_waiting_last_time;
  wire    [ 31: 0] ddr3_top_s1_readdata_from_sa_part_selected_by_negative_dbs;
  wire             empty_selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo;
  wire             full_selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo;
  wire             latency_load_value;
  wire             p1_pb_cpu_to_ddr3_top_m1_latency_counter;
  reg     [ 26: 0] pb_cpu_to_ddr3_top_m1_address_last_time;
  wire    [ 26: 0] pb_cpu_to_ddr3_top_m1_address_to_slave;
  reg              pb_cpu_to_ddr3_top_m1_burstcount_last_time;
  reg     [  3: 0] pb_cpu_to_ddr3_top_m1_byteenable_last_time;
  reg              pb_cpu_to_ddr3_top_m1_chipselect_last_time;
  wire             pb_cpu_to_ddr3_top_m1_is_granted_some_slave;
  reg              pb_cpu_to_ddr3_top_m1_latency_counter;
  reg              pb_cpu_to_ddr3_top_m1_read_but_no_slave_selected;
  reg              pb_cpu_to_ddr3_top_m1_read_last_time;
  wire    [ 31: 0] pb_cpu_to_ddr3_top_m1_readdata;
  wire             pb_cpu_to_ddr3_top_m1_readdatavalid;
  wire             pb_cpu_to_ddr3_top_m1_run;
  wire             pb_cpu_to_ddr3_top_m1_waitrequest;
  reg              pb_cpu_to_ddr3_top_m1_write_last_time;
  reg     [ 31: 0] pb_cpu_to_ddr3_top_m1_writedata_last_time;
  wire             pre_flush_pb_cpu_to_ddr3_top_m1_readdatavalid;
  wire             r_0;
  wire             read_selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo;
  wire             selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo_output;
  wire             selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo_output_ddr3_top_s1;
  wire             write_selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (pb_cpu_to_ddr3_top_m1_qualified_request_ddr3_top_s1 | ~pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1) & (pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1 | ~pb_cpu_to_ddr3_top_m1_qualified_request_ddr3_top_s1) & ((~pb_cpu_to_ddr3_top_m1_qualified_request_ddr3_top_s1 | ~pb_cpu_to_ddr3_top_m1_chipselect | (1 & ddr3_top_s1_waitrequest_n_from_sa & pb_cpu_to_ddr3_top_m1_chipselect))) & ((~pb_cpu_to_ddr3_top_m1_qualified_request_ddr3_top_s1 | ~pb_cpu_to_ddr3_top_m1_chipselect | (1 & ddr3_top_s1_waitrequest_n_from_sa & pb_cpu_to_ddr3_top_m1_chipselect)));

  //cascaded wait assignment, which is an e_assign
  assign pb_cpu_to_ddr3_top_m1_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign pb_cpu_to_ddr3_top_m1_address_to_slave = pb_cpu_to_ddr3_top_m1_address[26 : 0];

  //pb_cpu_to_ddr3_top_m1_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_ddr3_top_m1_read_but_no_slave_selected <= 0;
      else 
        pb_cpu_to_ddr3_top_m1_read_but_no_slave_selected <= (pb_cpu_to_ddr3_top_m1_read & pb_cpu_to_ddr3_top_m1_chipselect) & pb_cpu_to_ddr3_top_m1_run & ~pb_cpu_to_ddr3_top_m1_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign pb_cpu_to_ddr3_top_m1_is_granted_some_slave = pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_pb_cpu_to_ddr3_top_m1_readdatavalid = pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign pb_cpu_to_ddr3_top_m1_readdatavalid = pb_cpu_to_ddr3_top_m1_read_but_no_slave_selected |
    pre_flush_pb_cpu_to_ddr3_top_m1_readdatavalid;

  //Negative Dynamic Bus-sizing mux.
  //this mux selects the correct half of the 
  //wide data coming from the slave ddr3_top/s1 
  assign ddr3_top_s1_readdata_from_sa_part_selected_by_negative_dbs = ((selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo_output_ddr3_top_s1 == 0))? ddr3_top_s1_readdata_from_sa[31 : 0] :
    ddr3_top_s1_readdata_from_sa[63 : 32];

  //read_selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo fifo read, which is an e_mux
  assign read_selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo = pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1;

  //write_selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo fifo write, which is an e_mux
  assign write_selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo = (pb_cpu_to_ddr3_top_m1_read & pb_cpu_to_ddr3_top_m1_chipselect) & pb_cpu_to_ddr3_top_m1_run & pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1;

  assign selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo_output_ddr3_top_s1 = selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo_output;
  //selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo, which is an e_fifo_with_registered_outputs
  selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo_module selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (pb_cpu_to_ddr3_top_m1_address_to_slave[2]),
      .data_out             (selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo_output),
      .empty                (empty_selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo),
      .fifo_contains_ones_n (),
      .full                 (full_selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo),
      .read                 (read_selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (write_selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo)
    );

  //pb_cpu_to_ddr3_top/m1 readdata mux, which is an e_mux
  assign pb_cpu_to_ddr3_top_m1_readdata = ddr3_top_s1_readdata_from_sa_part_selected_by_negative_dbs;

  //actual waitrequest port, which is an e_assign
  assign pb_cpu_to_ddr3_top_m1_waitrequest = ~pb_cpu_to_ddr3_top_m1_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_ddr3_top_m1_latency_counter <= 0;
      else 
        pb_cpu_to_ddr3_top_m1_latency_counter <= p1_pb_cpu_to_ddr3_top_m1_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_pb_cpu_to_ddr3_top_m1_latency_counter = ((pb_cpu_to_ddr3_top_m1_run & (pb_cpu_to_ddr3_top_m1_read & pb_cpu_to_ddr3_top_m1_chipselect)))? latency_load_value :
    (pb_cpu_to_ddr3_top_m1_latency_counter)? pb_cpu_to_ddr3_top_m1_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pb_cpu_to_ddr3_top_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_ddr3_top_m1_address_last_time <= 0;
      else 
        pb_cpu_to_ddr3_top_m1_address_last_time <= pb_cpu_to_ddr3_top_m1_address;
    end


  //pb_cpu_to_ddr3_top/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= pb_cpu_to_ddr3_top_m1_waitrequest & pb_cpu_to_ddr3_top_m1_chipselect;
    end


  //pb_cpu_to_ddr3_top_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_ddr3_top_m1_address != pb_cpu_to_ddr3_top_m1_address_last_time))
        begin
          $write("%0d ns: pb_cpu_to_ddr3_top_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_ddr3_top_m1_chipselect check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_ddr3_top_m1_chipselect_last_time <= 0;
      else 
        pb_cpu_to_ddr3_top_m1_chipselect_last_time <= pb_cpu_to_ddr3_top_m1_chipselect;
    end


  //pb_cpu_to_ddr3_top_m1_chipselect matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_ddr3_top_m1_chipselect != pb_cpu_to_ddr3_top_m1_chipselect_last_time))
        begin
          $write("%0d ns: pb_cpu_to_ddr3_top_m1_chipselect did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_ddr3_top_m1_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_ddr3_top_m1_burstcount_last_time <= 0;
      else 
        pb_cpu_to_ddr3_top_m1_burstcount_last_time <= pb_cpu_to_ddr3_top_m1_burstcount;
    end


  //pb_cpu_to_ddr3_top_m1_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_ddr3_top_m1_burstcount != pb_cpu_to_ddr3_top_m1_burstcount_last_time))
        begin
          $write("%0d ns: pb_cpu_to_ddr3_top_m1_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_ddr3_top_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_ddr3_top_m1_byteenable_last_time <= 0;
      else 
        pb_cpu_to_ddr3_top_m1_byteenable_last_time <= pb_cpu_to_ddr3_top_m1_byteenable;
    end


  //pb_cpu_to_ddr3_top_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_ddr3_top_m1_byteenable != pb_cpu_to_ddr3_top_m1_byteenable_last_time))
        begin
          $write("%0d ns: pb_cpu_to_ddr3_top_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_ddr3_top_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_ddr3_top_m1_read_last_time <= 0;
      else 
        pb_cpu_to_ddr3_top_m1_read_last_time <= pb_cpu_to_ddr3_top_m1_read;
    end


  //pb_cpu_to_ddr3_top_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_ddr3_top_m1_read != pb_cpu_to_ddr3_top_m1_read_last_time))
        begin
          $write("%0d ns: pb_cpu_to_ddr3_top_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_ddr3_top_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_ddr3_top_m1_write_last_time <= 0;
      else 
        pb_cpu_to_ddr3_top_m1_write_last_time <= pb_cpu_to_ddr3_top_m1_write;
    end


  //pb_cpu_to_ddr3_top_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_ddr3_top_m1_write != pb_cpu_to_ddr3_top_m1_write_last_time))
        begin
          $write("%0d ns: pb_cpu_to_ddr3_top_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_ddr3_top_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_ddr3_top_m1_writedata_last_time <= 0;
      else 
        pb_cpu_to_ddr3_top_m1_writedata_last_time <= pb_cpu_to_ddr3_top_m1_writedata;
    end


  //pb_cpu_to_ddr3_top_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_ddr3_top_m1_writedata != pb_cpu_to_ddr3_top_m1_writedata_last_time) & (pb_cpu_to_ddr3_top_m1_write & pb_cpu_to_ddr3_top_m1_chipselect))
        begin
          $write("%0d ns: pb_cpu_to_ddr3_top_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end


  //selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo read when empty, which is an e_process
  always @(posedge clk)
    begin
      if (empty_selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo & read_selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo)
        begin
          $write("%0d ns: pb_cpu_to_ddr3_top/m1 negative rdv fifo selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo: read AND empty.\n", $time);
          $stop;
        end
    end


  //selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo write when full, which is an e_process
  always @(posedge clk)
    begin
      if (full_selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo & write_selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo & ~read_selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo)
        begin
          $write("%0d ns: pb_cpu_to_ddr3_top/m1 negative rdv fifo selecto_nrdv_pb_cpu_to_ddr3_top_m1_1_ddr3_top_s1_fifo: write AND full.\n", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pb_cpu_to_ddr3_top_bridge_arbitrator 
;



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_pb_cpu_to_fsm_s1_module (
                                                                 // inputs:
                                                                  clear_fifo,
                                                                  clk,
                                                                  data_in,
                                                                  read,
                                                                  reset_n,
                                                                  sync_reset,
                                                                  write,

                                                                 // outputs:
                                                                  data_out,
                                                                  empty,
                                                                  fifo_contains_ones_n,
                                                                  full
                                                               )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  wire             full_4;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_3;
  assign empty = !full_0;
  assign full_4 = 0;
  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    0;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_instruction_master_to_pb_cpu_to_fsm_s1_module (
                                                                        // inputs:
                                                                         clear_fifo,
                                                                         clk,
                                                                         data_in,
                                                                         read,
                                                                         reset_n,
                                                                         sync_reset,
                                                                         write,

                                                                        // outputs:
                                                                         data_out,
                                                                         empty,
                                                                         fifo_contains_ones_n,
                                                                         full
                                                                      )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  wire             full_4;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_3;
  assign empty = !full_0;
  assign full_4 = 0;
  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    0;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pb_cpu_to_fsm_s1_arbitrator (
                                     // inputs:
                                      clk,
                                      cpu_data_master_address_to_slave,
                                      cpu_data_master_byteenable,
                                      cpu_data_master_debugaccess,
                                      cpu_data_master_latency_counter,
                                      cpu_data_master_read,
                                      cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register,
                                      cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register,
                                      cpu_data_master_write,
                                      cpu_data_master_writedata,
                                      cpu_instruction_master_address_to_slave,
                                      cpu_instruction_master_latency_counter,
                                      cpu_instruction_master_read,
                                      cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register,
                                      pb_cpu_to_fsm_s1_endofpacket,
                                      pb_cpu_to_fsm_s1_readdata,
                                      pb_cpu_to_fsm_s1_readdatavalid,
                                      pb_cpu_to_fsm_s1_waitrequest,
                                      reset_n,

                                     // outputs:
                                      cpu_data_master_granted_pb_cpu_to_fsm_s1,
                                      cpu_data_master_qualified_request_pb_cpu_to_fsm_s1,
                                      cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1,
                                      cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register,
                                      cpu_data_master_requests_pb_cpu_to_fsm_s1,
                                      cpu_instruction_master_granted_pb_cpu_to_fsm_s1,
                                      cpu_instruction_master_qualified_request_pb_cpu_to_fsm_s1,
                                      cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1,
                                      cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register,
                                      cpu_instruction_master_requests_pb_cpu_to_fsm_s1,
                                      d1_pb_cpu_to_fsm_s1_end_xfer,
                                      pb_cpu_to_fsm_s1_address,
                                      pb_cpu_to_fsm_s1_arbiterlock,
                                      pb_cpu_to_fsm_s1_arbiterlock2,
                                      pb_cpu_to_fsm_s1_burstcount,
                                      pb_cpu_to_fsm_s1_byteenable,
                                      pb_cpu_to_fsm_s1_chipselect,
                                      pb_cpu_to_fsm_s1_debugaccess,
                                      pb_cpu_to_fsm_s1_endofpacket_from_sa,
                                      pb_cpu_to_fsm_s1_nativeaddress,
                                      pb_cpu_to_fsm_s1_read,
                                      pb_cpu_to_fsm_s1_readdata_from_sa,
                                      pb_cpu_to_fsm_s1_reset_n,
                                      pb_cpu_to_fsm_s1_waitrequest_from_sa,
                                      pb_cpu_to_fsm_s1_write,
                                      pb_cpu_to_fsm_s1_writedata
                                   )
;

  output           cpu_data_master_granted_pb_cpu_to_fsm_s1;
  output           cpu_data_master_qualified_request_pb_cpu_to_fsm_s1;
  output           cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1;
  output           cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register;
  output           cpu_data_master_requests_pb_cpu_to_fsm_s1;
  output           cpu_instruction_master_granted_pb_cpu_to_fsm_s1;
  output           cpu_instruction_master_qualified_request_pb_cpu_to_fsm_s1;
  output           cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1;
  output           cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register;
  output           cpu_instruction_master_requests_pb_cpu_to_fsm_s1;
  output           d1_pb_cpu_to_fsm_s1_end_xfer;
  output  [ 23: 0] pb_cpu_to_fsm_s1_address;
  output           pb_cpu_to_fsm_s1_arbiterlock;
  output           pb_cpu_to_fsm_s1_arbiterlock2;
  output           pb_cpu_to_fsm_s1_burstcount;
  output  [  3: 0] pb_cpu_to_fsm_s1_byteenable;
  output           pb_cpu_to_fsm_s1_chipselect;
  output           pb_cpu_to_fsm_s1_debugaccess;
  output           pb_cpu_to_fsm_s1_endofpacket_from_sa;
  output  [ 23: 0] pb_cpu_to_fsm_s1_nativeaddress;
  output           pb_cpu_to_fsm_s1_read;
  output  [ 31: 0] pb_cpu_to_fsm_s1_readdata_from_sa;
  output           pb_cpu_to_fsm_s1_reset_n;
  output           pb_cpu_to_fsm_s1_waitrequest_from_sa;
  output           pb_cpu_to_fsm_s1_write;
  output  [ 31: 0] pb_cpu_to_fsm_s1_writedata;
  input            clk;
  input   [ 28: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register;
  input            cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 28: 0] cpu_instruction_master_address_to_slave;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register;
  input            pb_cpu_to_fsm_s1_endofpacket;
  input   [ 31: 0] pb_cpu_to_fsm_s1_readdata;
  input            pb_cpu_to_fsm_s1_readdatavalid;
  input            pb_cpu_to_fsm_s1_waitrequest;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_pb_cpu_to_fsm_s1;
  wire             cpu_data_master_qualified_request_pb_cpu_to_fsm_s1;
  wire             cpu_data_master_rdv_fifo_empty_pb_cpu_to_fsm_s1;
  wire             cpu_data_master_rdv_fifo_output_from_pb_cpu_to_fsm_s1;
  wire             cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1;
  wire             cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register;
  wire             cpu_data_master_requests_pb_cpu_to_fsm_s1;
  wire             cpu_data_master_saved_grant_pb_cpu_to_fsm_s1;
  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_pb_cpu_to_fsm_s1;
  wire             cpu_instruction_master_qualified_request_pb_cpu_to_fsm_s1;
  wire             cpu_instruction_master_rdv_fifo_empty_pb_cpu_to_fsm_s1;
  wire             cpu_instruction_master_rdv_fifo_output_from_pb_cpu_to_fsm_s1;
  wire             cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1;
  wire             cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register;
  wire             cpu_instruction_master_requests_pb_cpu_to_fsm_s1;
  wire             cpu_instruction_master_saved_grant_pb_cpu_to_fsm_s1;
  reg              d1_pb_cpu_to_fsm_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_pb_cpu_to_fsm_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_data_master_granted_slave_pb_cpu_to_fsm_s1;
  reg              last_cycle_cpu_instruction_master_granted_slave_pb_cpu_to_fsm_s1;
  wire    [ 23: 0] pb_cpu_to_fsm_s1_address;
  wire             pb_cpu_to_fsm_s1_allgrants;
  wire             pb_cpu_to_fsm_s1_allow_new_arb_cycle;
  wire             pb_cpu_to_fsm_s1_any_bursting_master_saved_grant;
  wire             pb_cpu_to_fsm_s1_any_continuerequest;
  reg     [  1: 0] pb_cpu_to_fsm_s1_arb_addend;
  wire             pb_cpu_to_fsm_s1_arb_counter_enable;
  reg     [  3: 0] pb_cpu_to_fsm_s1_arb_share_counter;
  wire    [  3: 0] pb_cpu_to_fsm_s1_arb_share_counter_next_value;
  wire    [  3: 0] pb_cpu_to_fsm_s1_arb_share_set_values;
  wire    [  1: 0] pb_cpu_to_fsm_s1_arb_winner;
  wire             pb_cpu_to_fsm_s1_arbiterlock;
  wire             pb_cpu_to_fsm_s1_arbiterlock2;
  wire             pb_cpu_to_fsm_s1_arbitration_holdoff_internal;
  wire             pb_cpu_to_fsm_s1_beginbursttransfer_internal;
  wire             pb_cpu_to_fsm_s1_begins_xfer;
  wire             pb_cpu_to_fsm_s1_burstcount;
  wire    [  3: 0] pb_cpu_to_fsm_s1_byteenable;
  wire             pb_cpu_to_fsm_s1_chipselect;
  wire    [  3: 0] pb_cpu_to_fsm_s1_chosen_master_double_vector;
  wire    [  1: 0] pb_cpu_to_fsm_s1_chosen_master_rot_left;
  wire             pb_cpu_to_fsm_s1_debugaccess;
  wire             pb_cpu_to_fsm_s1_end_xfer;
  wire             pb_cpu_to_fsm_s1_endofpacket_from_sa;
  wire             pb_cpu_to_fsm_s1_firsttransfer;
  wire    [  1: 0] pb_cpu_to_fsm_s1_grant_vector;
  wire             pb_cpu_to_fsm_s1_in_a_read_cycle;
  wire             pb_cpu_to_fsm_s1_in_a_write_cycle;
  wire    [  1: 0] pb_cpu_to_fsm_s1_master_qreq_vector;
  wire             pb_cpu_to_fsm_s1_move_on_to_next_transaction;
  wire    [ 23: 0] pb_cpu_to_fsm_s1_nativeaddress;
  wire             pb_cpu_to_fsm_s1_non_bursting_master_requests;
  wire             pb_cpu_to_fsm_s1_read;
  wire    [ 31: 0] pb_cpu_to_fsm_s1_readdata_from_sa;
  wire             pb_cpu_to_fsm_s1_readdatavalid_from_sa;
  reg              pb_cpu_to_fsm_s1_reg_firsttransfer;
  wire             pb_cpu_to_fsm_s1_reset_n;
  reg     [  1: 0] pb_cpu_to_fsm_s1_saved_chosen_master_vector;
  reg              pb_cpu_to_fsm_s1_slavearbiterlockenable;
  wire             pb_cpu_to_fsm_s1_slavearbiterlockenable2;
  wire             pb_cpu_to_fsm_s1_unreg_firsttransfer;
  wire             pb_cpu_to_fsm_s1_waitrequest_from_sa;
  wire             pb_cpu_to_fsm_s1_waits_for_read;
  wire             pb_cpu_to_fsm_s1_waits_for_write;
  wire             pb_cpu_to_fsm_s1_write;
  wire    [ 31: 0] pb_cpu_to_fsm_s1_writedata;
  wire    [ 28: 0] shifted_address_to_pb_cpu_to_fsm_s1_from_cpu_data_master;
  wire    [ 28: 0] shifted_address_to_pb_cpu_to_fsm_s1_from_cpu_instruction_master;
  wire             wait_for_pb_cpu_to_fsm_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~pb_cpu_to_fsm_s1_end_xfer;
    end


  assign pb_cpu_to_fsm_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_pb_cpu_to_fsm_s1 | cpu_instruction_master_qualified_request_pb_cpu_to_fsm_s1));
  //assign pb_cpu_to_fsm_s1_readdatavalid_from_sa = pb_cpu_to_fsm_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_cpu_to_fsm_s1_readdatavalid_from_sa = pb_cpu_to_fsm_s1_readdatavalid;

  //assign pb_cpu_to_fsm_s1_readdata_from_sa = pb_cpu_to_fsm_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_cpu_to_fsm_s1_readdata_from_sa = pb_cpu_to_fsm_s1_readdata;

  assign cpu_data_master_requests_pb_cpu_to_fsm_s1 = ({cpu_data_master_address_to_slave[28 : 26] , 26'b0} == 29'h0) & (cpu_data_master_read | cpu_data_master_write);
  //assign pb_cpu_to_fsm_s1_waitrequest_from_sa = pb_cpu_to_fsm_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_cpu_to_fsm_s1_waitrequest_from_sa = pb_cpu_to_fsm_s1_waitrequest;

  //pb_cpu_to_fsm_s1_arb_share_counter set values, which is an e_mux
  assign pb_cpu_to_fsm_s1_arb_share_set_values = (cpu_data_master_granted_pb_cpu_to_fsm_s1)? 8 :
    (cpu_instruction_master_granted_pb_cpu_to_fsm_s1)? 8 :
    (cpu_data_master_granted_pb_cpu_to_fsm_s1)? 8 :
    (cpu_instruction_master_granted_pb_cpu_to_fsm_s1)? 8 :
    (cpu_data_master_granted_pb_cpu_to_fsm_s1)? 8 :
    (cpu_instruction_master_granted_pb_cpu_to_fsm_s1)? 8 :
    1;

  //pb_cpu_to_fsm_s1_non_bursting_master_requests mux, which is an e_mux
  assign pb_cpu_to_fsm_s1_non_bursting_master_requests = cpu_data_master_requests_pb_cpu_to_fsm_s1 |
    cpu_instruction_master_requests_pb_cpu_to_fsm_s1 |
    cpu_data_master_requests_pb_cpu_to_fsm_s1 |
    cpu_instruction_master_requests_pb_cpu_to_fsm_s1 |
    cpu_data_master_requests_pb_cpu_to_fsm_s1 |
    cpu_instruction_master_requests_pb_cpu_to_fsm_s1;

  //pb_cpu_to_fsm_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign pb_cpu_to_fsm_s1_any_bursting_master_saved_grant = 0;

  //pb_cpu_to_fsm_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign pb_cpu_to_fsm_s1_arb_share_counter_next_value = pb_cpu_to_fsm_s1_firsttransfer ? (pb_cpu_to_fsm_s1_arb_share_set_values - 1) : |pb_cpu_to_fsm_s1_arb_share_counter ? (pb_cpu_to_fsm_s1_arb_share_counter - 1) : 0;

  //pb_cpu_to_fsm_s1_allgrants all slave grants, which is an e_mux
  assign pb_cpu_to_fsm_s1_allgrants = (|pb_cpu_to_fsm_s1_grant_vector) |
    (|pb_cpu_to_fsm_s1_grant_vector) |
    (|pb_cpu_to_fsm_s1_grant_vector) |
    (|pb_cpu_to_fsm_s1_grant_vector) |
    (|pb_cpu_to_fsm_s1_grant_vector) |
    (|pb_cpu_to_fsm_s1_grant_vector);

  //pb_cpu_to_fsm_s1_end_xfer assignment, which is an e_assign
  assign pb_cpu_to_fsm_s1_end_xfer = ~(pb_cpu_to_fsm_s1_waits_for_read | pb_cpu_to_fsm_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_pb_cpu_to_fsm_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_pb_cpu_to_fsm_s1 = pb_cpu_to_fsm_s1_end_xfer & (~pb_cpu_to_fsm_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //pb_cpu_to_fsm_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign pb_cpu_to_fsm_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_pb_cpu_to_fsm_s1 & pb_cpu_to_fsm_s1_allgrants) | (end_xfer_arb_share_counter_term_pb_cpu_to_fsm_s1 & ~pb_cpu_to_fsm_s1_non_bursting_master_requests);

  //pb_cpu_to_fsm_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_s1_arb_share_counter <= 0;
      else if (pb_cpu_to_fsm_s1_arb_counter_enable)
          pb_cpu_to_fsm_s1_arb_share_counter <= pb_cpu_to_fsm_s1_arb_share_counter_next_value;
    end


  //pb_cpu_to_fsm_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_s1_slavearbiterlockenable <= 0;
      else if ((|pb_cpu_to_fsm_s1_master_qreq_vector & end_xfer_arb_share_counter_term_pb_cpu_to_fsm_s1) | (end_xfer_arb_share_counter_term_pb_cpu_to_fsm_s1 & ~pb_cpu_to_fsm_s1_non_bursting_master_requests))
          pb_cpu_to_fsm_s1_slavearbiterlockenable <= |pb_cpu_to_fsm_s1_arb_share_counter_next_value;
    end


  //cpu/data_master pb_cpu_to_fsm/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = pb_cpu_to_fsm_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //pb_cpu_to_fsm_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign pb_cpu_to_fsm_s1_slavearbiterlockenable2 = |pb_cpu_to_fsm_s1_arb_share_counter_next_value;

  //cpu/data_master pb_cpu_to_fsm/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = pb_cpu_to_fsm_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //cpu/instruction_master pb_cpu_to_fsm/s1 arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = pb_cpu_to_fsm_s1_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //cpu/instruction_master pb_cpu_to_fsm/s1 arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = pb_cpu_to_fsm_s1_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //cpu/instruction_master granted pb_cpu_to_fsm/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_instruction_master_granted_slave_pb_cpu_to_fsm_s1 <= 0;
      else 
        last_cycle_cpu_instruction_master_granted_slave_pb_cpu_to_fsm_s1 <= cpu_instruction_master_saved_grant_pb_cpu_to_fsm_s1 ? 1 : (pb_cpu_to_fsm_s1_arbitration_holdoff_internal | ~cpu_instruction_master_requests_pb_cpu_to_fsm_s1) ? 0 : last_cycle_cpu_instruction_master_granted_slave_pb_cpu_to_fsm_s1;
    end


  //cpu_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_instruction_master_continuerequest = last_cycle_cpu_instruction_master_granted_slave_pb_cpu_to_fsm_s1 & cpu_instruction_master_requests_pb_cpu_to_fsm_s1;

  //pb_cpu_to_fsm_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign pb_cpu_to_fsm_s1_any_continuerequest = cpu_instruction_master_continuerequest |
    cpu_data_master_continuerequest;

  assign cpu_data_master_qualified_request_pb_cpu_to_fsm_s1 = cpu_data_master_requests_pb_cpu_to_fsm_s1 & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register) | (|cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register))) | cpu_instruction_master_arbiterlock);
  //unique name for pb_cpu_to_fsm_s1_move_on_to_next_transaction, which is an e_assign
  assign pb_cpu_to_fsm_s1_move_on_to_next_transaction = pb_cpu_to_fsm_s1_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_pb_cpu_to_fsm_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_pb_cpu_to_fsm_s1_module rdv_fifo_for_cpu_data_master_to_pb_cpu_to_fsm_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_pb_cpu_to_fsm_s1),
      .data_out             (cpu_data_master_rdv_fifo_output_from_pb_cpu_to_fsm_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_pb_cpu_to_fsm_s1),
      .full                 (),
      .read                 (pb_cpu_to_fsm_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~pb_cpu_to_fsm_s1_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register = ~cpu_data_master_rdv_fifo_empty_pb_cpu_to_fsm_s1;
  //local readdatavalid cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1 = (pb_cpu_to_fsm_s1_readdatavalid_from_sa & cpu_data_master_rdv_fifo_output_from_pb_cpu_to_fsm_s1) & ~ cpu_data_master_rdv_fifo_empty_pb_cpu_to_fsm_s1;

  //pb_cpu_to_fsm_s1_writedata mux, which is an e_mux
  assign pb_cpu_to_fsm_s1_writedata = cpu_data_master_writedata;

  //assign pb_cpu_to_fsm_s1_endofpacket_from_sa = pb_cpu_to_fsm_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_cpu_to_fsm_s1_endofpacket_from_sa = pb_cpu_to_fsm_s1_endofpacket;

  assign cpu_instruction_master_requests_pb_cpu_to_fsm_s1 = (({cpu_instruction_master_address_to_slave[28 : 26] , 26'b0} == 29'h0) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //cpu/data_master granted pb_cpu_to_fsm/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_data_master_granted_slave_pb_cpu_to_fsm_s1 <= 0;
      else 
        last_cycle_cpu_data_master_granted_slave_pb_cpu_to_fsm_s1 <= cpu_data_master_saved_grant_pb_cpu_to_fsm_s1 ? 1 : (pb_cpu_to_fsm_s1_arbitration_holdoff_internal | ~cpu_data_master_requests_pb_cpu_to_fsm_s1) ? 0 : last_cycle_cpu_data_master_granted_slave_pb_cpu_to_fsm_s1;
    end


  //cpu_data_master_continuerequest continued request, which is an e_mux
  assign cpu_data_master_continuerequest = last_cycle_cpu_data_master_granted_slave_pb_cpu_to_fsm_s1 & cpu_data_master_requests_pb_cpu_to_fsm_s1;

  assign cpu_instruction_master_qualified_request_pb_cpu_to_fsm_s1 = cpu_instruction_master_requests_pb_cpu_to_fsm_s1 & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (1 < cpu_instruction_master_latency_counter) | (|cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register))) | cpu_data_master_arbiterlock);
  //rdv_fifo_for_cpu_instruction_master_to_pb_cpu_to_fsm_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_pb_cpu_to_fsm_s1_module rdv_fifo_for_cpu_instruction_master_to_pb_cpu_to_fsm_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_instruction_master_granted_pb_cpu_to_fsm_s1),
      .data_out             (cpu_instruction_master_rdv_fifo_output_from_pb_cpu_to_fsm_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_instruction_master_rdv_fifo_empty_pb_cpu_to_fsm_s1),
      .full                 (),
      .read                 (pb_cpu_to_fsm_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~pb_cpu_to_fsm_s1_waits_for_read)
    );

  assign cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register = ~cpu_instruction_master_rdv_fifo_empty_pb_cpu_to_fsm_s1;
  //local readdatavalid cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1, which is an e_mux
  assign cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1 = (pb_cpu_to_fsm_s1_readdatavalid_from_sa & cpu_instruction_master_rdv_fifo_output_from_pb_cpu_to_fsm_s1) & ~ cpu_instruction_master_rdv_fifo_empty_pb_cpu_to_fsm_s1;

  //allow new arb cycle for pb_cpu_to_fsm/s1, which is an e_assign
  assign pb_cpu_to_fsm_s1_allow_new_arb_cycle = ~cpu_data_master_arbiterlock & ~cpu_instruction_master_arbiterlock;

  //cpu/instruction_master assignment into master qualified-requests vector for pb_cpu_to_fsm/s1, which is an e_assign
  assign pb_cpu_to_fsm_s1_master_qreq_vector[0] = cpu_instruction_master_qualified_request_pb_cpu_to_fsm_s1;

  //cpu/instruction_master grant pb_cpu_to_fsm/s1, which is an e_assign
  assign cpu_instruction_master_granted_pb_cpu_to_fsm_s1 = pb_cpu_to_fsm_s1_grant_vector[0];

  //cpu/instruction_master saved-grant pb_cpu_to_fsm/s1, which is an e_assign
  assign cpu_instruction_master_saved_grant_pb_cpu_to_fsm_s1 = pb_cpu_to_fsm_s1_arb_winner[0] && cpu_instruction_master_requests_pb_cpu_to_fsm_s1;

  //cpu/data_master assignment into master qualified-requests vector for pb_cpu_to_fsm/s1, which is an e_assign
  assign pb_cpu_to_fsm_s1_master_qreq_vector[1] = cpu_data_master_qualified_request_pb_cpu_to_fsm_s1;

  //cpu/data_master grant pb_cpu_to_fsm/s1, which is an e_assign
  assign cpu_data_master_granted_pb_cpu_to_fsm_s1 = pb_cpu_to_fsm_s1_grant_vector[1];

  //cpu/data_master saved-grant pb_cpu_to_fsm/s1, which is an e_assign
  assign cpu_data_master_saved_grant_pb_cpu_to_fsm_s1 = pb_cpu_to_fsm_s1_arb_winner[1] && cpu_data_master_requests_pb_cpu_to_fsm_s1;

  //pb_cpu_to_fsm/s1 chosen-master double-vector, which is an e_assign
  assign pb_cpu_to_fsm_s1_chosen_master_double_vector = {pb_cpu_to_fsm_s1_master_qreq_vector, pb_cpu_to_fsm_s1_master_qreq_vector} & ({~pb_cpu_to_fsm_s1_master_qreq_vector, ~pb_cpu_to_fsm_s1_master_qreq_vector} + pb_cpu_to_fsm_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign pb_cpu_to_fsm_s1_arb_winner = (pb_cpu_to_fsm_s1_allow_new_arb_cycle & | pb_cpu_to_fsm_s1_grant_vector) ? pb_cpu_to_fsm_s1_grant_vector : pb_cpu_to_fsm_s1_saved_chosen_master_vector;

  //saved pb_cpu_to_fsm_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_s1_saved_chosen_master_vector <= 0;
      else if (pb_cpu_to_fsm_s1_allow_new_arb_cycle)
          pb_cpu_to_fsm_s1_saved_chosen_master_vector <= |pb_cpu_to_fsm_s1_grant_vector ? pb_cpu_to_fsm_s1_grant_vector : pb_cpu_to_fsm_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign pb_cpu_to_fsm_s1_grant_vector = {(pb_cpu_to_fsm_s1_chosen_master_double_vector[1] | pb_cpu_to_fsm_s1_chosen_master_double_vector[3]),
    (pb_cpu_to_fsm_s1_chosen_master_double_vector[0] | pb_cpu_to_fsm_s1_chosen_master_double_vector[2])};

  //pb_cpu_to_fsm/s1 chosen master rotated left, which is an e_assign
  assign pb_cpu_to_fsm_s1_chosen_master_rot_left = (pb_cpu_to_fsm_s1_arb_winner << 1) ? (pb_cpu_to_fsm_s1_arb_winner << 1) : 1;

  //pb_cpu_to_fsm/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_s1_arb_addend <= 1;
      else if (|pb_cpu_to_fsm_s1_grant_vector)
          pb_cpu_to_fsm_s1_arb_addend <= pb_cpu_to_fsm_s1_end_xfer? pb_cpu_to_fsm_s1_chosen_master_rot_left : pb_cpu_to_fsm_s1_grant_vector;
    end


  //pb_cpu_to_fsm_s1_reset_n assignment, which is an e_assign
  assign pb_cpu_to_fsm_s1_reset_n = reset_n;

  assign pb_cpu_to_fsm_s1_chipselect = cpu_data_master_granted_pb_cpu_to_fsm_s1 | cpu_instruction_master_granted_pb_cpu_to_fsm_s1;
  //pb_cpu_to_fsm_s1_firsttransfer first transaction, which is an e_assign
  assign pb_cpu_to_fsm_s1_firsttransfer = pb_cpu_to_fsm_s1_begins_xfer ? pb_cpu_to_fsm_s1_unreg_firsttransfer : pb_cpu_to_fsm_s1_reg_firsttransfer;

  //pb_cpu_to_fsm_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign pb_cpu_to_fsm_s1_unreg_firsttransfer = ~(pb_cpu_to_fsm_s1_slavearbiterlockenable & pb_cpu_to_fsm_s1_any_continuerequest);

  //pb_cpu_to_fsm_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_s1_reg_firsttransfer <= 1'b1;
      else if (pb_cpu_to_fsm_s1_begins_xfer)
          pb_cpu_to_fsm_s1_reg_firsttransfer <= pb_cpu_to_fsm_s1_unreg_firsttransfer;
    end


  //pb_cpu_to_fsm_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign pb_cpu_to_fsm_s1_beginbursttransfer_internal = pb_cpu_to_fsm_s1_begins_xfer;

  //pb_cpu_to_fsm_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign pb_cpu_to_fsm_s1_arbitration_holdoff_internal = pb_cpu_to_fsm_s1_begins_xfer & pb_cpu_to_fsm_s1_firsttransfer;

  //pb_cpu_to_fsm_s1_read assignment, which is an e_mux
  assign pb_cpu_to_fsm_s1_read = (cpu_data_master_granted_pb_cpu_to_fsm_s1 & cpu_data_master_read) | (cpu_instruction_master_granted_pb_cpu_to_fsm_s1 & cpu_instruction_master_read);

  //pb_cpu_to_fsm_s1_write assignment, which is an e_mux
  assign pb_cpu_to_fsm_s1_write = cpu_data_master_granted_pb_cpu_to_fsm_s1 & cpu_data_master_write;

  assign shifted_address_to_pb_cpu_to_fsm_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //pb_cpu_to_fsm_s1_address mux, which is an e_mux
  assign pb_cpu_to_fsm_s1_address = (cpu_data_master_granted_pb_cpu_to_fsm_s1)? (shifted_address_to_pb_cpu_to_fsm_s1_from_cpu_data_master >> 2) :
    (shifted_address_to_pb_cpu_to_fsm_s1_from_cpu_instruction_master >> 2);

  assign shifted_address_to_pb_cpu_to_fsm_s1_from_cpu_instruction_master = cpu_instruction_master_address_to_slave;
  //slaveid pb_cpu_to_fsm_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign pb_cpu_to_fsm_s1_nativeaddress = (cpu_data_master_granted_pb_cpu_to_fsm_s1)? (cpu_data_master_address_to_slave >> 2) :
    (cpu_instruction_master_address_to_slave >> 2);

  //d1_pb_cpu_to_fsm_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_pb_cpu_to_fsm_s1_end_xfer <= 1;
      else 
        d1_pb_cpu_to_fsm_s1_end_xfer <= pb_cpu_to_fsm_s1_end_xfer;
    end


  //pb_cpu_to_fsm_s1_waits_for_read in a cycle, which is an e_mux
  assign pb_cpu_to_fsm_s1_waits_for_read = pb_cpu_to_fsm_s1_in_a_read_cycle & pb_cpu_to_fsm_s1_waitrequest_from_sa;

  //pb_cpu_to_fsm_s1_in_a_read_cycle assignment, which is an e_assign
  assign pb_cpu_to_fsm_s1_in_a_read_cycle = (cpu_data_master_granted_pb_cpu_to_fsm_s1 & cpu_data_master_read) | (cpu_instruction_master_granted_pb_cpu_to_fsm_s1 & cpu_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = pb_cpu_to_fsm_s1_in_a_read_cycle;

  //pb_cpu_to_fsm_s1_waits_for_write in a cycle, which is an e_mux
  assign pb_cpu_to_fsm_s1_waits_for_write = pb_cpu_to_fsm_s1_in_a_write_cycle & pb_cpu_to_fsm_s1_waitrequest_from_sa;

  //pb_cpu_to_fsm_s1_in_a_write_cycle assignment, which is an e_assign
  assign pb_cpu_to_fsm_s1_in_a_write_cycle = cpu_data_master_granted_pb_cpu_to_fsm_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = pb_cpu_to_fsm_s1_in_a_write_cycle;

  assign wait_for_pb_cpu_to_fsm_s1_counter = 0;
  //pb_cpu_to_fsm_s1_byteenable byte enable port mux, which is an e_mux
  assign pb_cpu_to_fsm_s1_byteenable = (cpu_data_master_granted_pb_cpu_to_fsm_s1)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign pb_cpu_to_fsm_s1_burstcount = 1;

  //pb_cpu_to_fsm/s1 arbiterlock assigned from _handle_arbiterlock, which is an e_mux
  assign pb_cpu_to_fsm_s1_arbiterlock = (cpu_data_master_arbiterlock)? cpu_data_master_arbiterlock :
    cpu_instruction_master_arbiterlock;

  //pb_cpu_to_fsm/s1 arbiterlock2 assigned from _handle_arbiterlock2, which is an e_mux
  assign pb_cpu_to_fsm_s1_arbiterlock2 = (cpu_data_master_arbiterlock2)? cpu_data_master_arbiterlock2 :
    cpu_instruction_master_arbiterlock2;

  //debugaccess mux, which is an e_mux
  assign pb_cpu_to_fsm_s1_debugaccess = (cpu_data_master_granted_pb_cpu_to_fsm_s1)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pb_cpu_to_fsm/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_granted_pb_cpu_to_fsm_s1 + cpu_instruction_master_granted_pb_cpu_to_fsm_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_saved_grant_pb_cpu_to_fsm_s1 + cpu_instruction_master_saved_grant_pb_cpu_to_fsm_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pb_cpu_to_fsm_m1_arbitrator (
                                     // inputs:
                                      clk,
                                      d1_tb_fsm_avalon_slave_end_xfer,
                                      ext_flash_1_s1_wait_counter_eq_0,
                                      ext_flash_s1_wait_counter_eq_0,
                                      incoming_tb_fsm_data_with_Xs_converted_to_0,
                                      pb_cpu_to_fsm_m1_address,
                                      pb_cpu_to_fsm_m1_burstcount,
                                      pb_cpu_to_fsm_m1_byteenable,
                                      pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1,
                                      pb_cpu_to_fsm_m1_byteenable_ext_flash_s1,
                                      pb_cpu_to_fsm_m1_chipselect,
                                      pb_cpu_to_fsm_m1_granted_ext_flash_1_s1,
                                      pb_cpu_to_fsm_m1_granted_ext_flash_s1,
                                      pb_cpu_to_fsm_m1_qualified_request_ext_flash_1_s1,
                                      pb_cpu_to_fsm_m1_qualified_request_ext_flash_s1,
                                      pb_cpu_to_fsm_m1_read,
                                      pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1,
                                      pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1,
                                      pb_cpu_to_fsm_m1_requests_ext_flash_1_s1,
                                      pb_cpu_to_fsm_m1_requests_ext_flash_s1,
                                      pb_cpu_to_fsm_m1_write,
                                      pb_cpu_to_fsm_m1_writedata,
                                      reset_n,

                                     // outputs:
                                      pb_cpu_to_fsm_m1_address_to_slave,
                                      pb_cpu_to_fsm_m1_dbs_address,
                                      pb_cpu_to_fsm_m1_dbs_write_16,
                                      pb_cpu_to_fsm_m1_latency_counter,
                                      pb_cpu_to_fsm_m1_readdata,
                                      pb_cpu_to_fsm_m1_readdatavalid,
                                      pb_cpu_to_fsm_m1_waitrequest
                                   )
;

  output  [ 25: 0] pb_cpu_to_fsm_m1_address_to_slave;
  output  [  1: 0] pb_cpu_to_fsm_m1_dbs_address;
  output  [ 15: 0] pb_cpu_to_fsm_m1_dbs_write_16;
  output  [  1: 0] pb_cpu_to_fsm_m1_latency_counter;
  output  [ 31: 0] pb_cpu_to_fsm_m1_readdata;
  output           pb_cpu_to_fsm_m1_readdatavalid;
  output           pb_cpu_to_fsm_m1_waitrequest;
  input            clk;
  input            d1_tb_fsm_avalon_slave_end_xfer;
  input            ext_flash_1_s1_wait_counter_eq_0;
  input            ext_flash_s1_wait_counter_eq_0;
  input   [ 15: 0] incoming_tb_fsm_data_with_Xs_converted_to_0;
  input   [ 25: 0] pb_cpu_to_fsm_m1_address;
  input            pb_cpu_to_fsm_m1_burstcount;
  input   [  3: 0] pb_cpu_to_fsm_m1_byteenable;
  input   [  1: 0] pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1;
  input   [  1: 0] pb_cpu_to_fsm_m1_byteenable_ext_flash_s1;
  input            pb_cpu_to_fsm_m1_chipselect;
  input            pb_cpu_to_fsm_m1_granted_ext_flash_1_s1;
  input            pb_cpu_to_fsm_m1_granted_ext_flash_s1;
  input            pb_cpu_to_fsm_m1_qualified_request_ext_flash_1_s1;
  input            pb_cpu_to_fsm_m1_qualified_request_ext_flash_s1;
  input            pb_cpu_to_fsm_m1_read;
  input            pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1;
  input            pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1;
  input            pb_cpu_to_fsm_m1_requests_ext_flash_1_s1;
  input            pb_cpu_to_fsm_m1_requests_ext_flash_s1;
  input            pb_cpu_to_fsm_m1_write;
  input   [ 31: 0] pb_cpu_to_fsm_m1_writedata;
  input            reset_n;

  reg              active_and_waiting_last_time;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [ 15: 0] dbs_latent_16_reg_segment_0;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  wire    [  1: 0] latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_0;
  wire    [  1: 0] p1_pb_cpu_to_fsm_m1_latency_counter;
  reg     [ 25: 0] pb_cpu_to_fsm_m1_address_last_time;
  wire    [ 25: 0] pb_cpu_to_fsm_m1_address_to_slave;
  reg              pb_cpu_to_fsm_m1_burstcount_last_time;
  reg     [  3: 0] pb_cpu_to_fsm_m1_byteenable_last_time;
  reg              pb_cpu_to_fsm_m1_chipselect_last_time;
  reg     [  1: 0] pb_cpu_to_fsm_m1_dbs_address;
  wire    [  1: 0] pb_cpu_to_fsm_m1_dbs_increment;
  reg     [  1: 0] pb_cpu_to_fsm_m1_dbs_rdv_counter;
  wire    [  1: 0] pb_cpu_to_fsm_m1_dbs_rdv_counter_inc;
  wire    [ 15: 0] pb_cpu_to_fsm_m1_dbs_write_16;
  wire             pb_cpu_to_fsm_m1_is_granted_some_slave;
  reg     [  1: 0] pb_cpu_to_fsm_m1_latency_counter;
  wire    [  1: 0] pb_cpu_to_fsm_m1_next_dbs_rdv_counter;
  reg              pb_cpu_to_fsm_m1_read_but_no_slave_selected;
  reg              pb_cpu_to_fsm_m1_read_last_time;
  wire    [ 31: 0] pb_cpu_to_fsm_m1_readdata;
  wire             pb_cpu_to_fsm_m1_readdatavalid;
  wire             pb_cpu_to_fsm_m1_run;
  wire             pb_cpu_to_fsm_m1_waitrequest;
  reg              pb_cpu_to_fsm_m1_write_last_time;
  reg     [ 31: 0] pb_cpu_to_fsm_m1_writedata_last_time;
  wire             pre_dbs_count_enable;
  wire             pre_flush_pb_cpu_to_fsm_m1_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & ((pb_cpu_to_fsm_m1_qualified_request_ext_flash_1_s1 | ((pb_cpu_to_fsm_m1_write & pb_cpu_to_fsm_m1_chipselect) & !pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1 & pb_cpu_to_fsm_m1_dbs_address[1]) | ~pb_cpu_to_fsm_m1_requests_ext_flash_1_s1)) & ((pb_cpu_to_fsm_m1_qualified_request_ext_flash_s1 | ((pb_cpu_to_fsm_m1_write & pb_cpu_to_fsm_m1_chipselect) & !pb_cpu_to_fsm_m1_byteenable_ext_flash_s1 & pb_cpu_to_fsm_m1_dbs_address[1]) | ~pb_cpu_to_fsm_m1_requests_ext_flash_s1)) & ((~pb_cpu_to_fsm_m1_qualified_request_ext_flash_1_s1 | ~(pb_cpu_to_fsm_m1_read & pb_cpu_to_fsm_m1_chipselect) | (1 & ((ext_flash_1_s1_wait_counter_eq_0 & ~d1_tb_fsm_avalon_slave_end_xfer)) & (pb_cpu_to_fsm_m1_dbs_address[1]) & (pb_cpu_to_fsm_m1_read & pb_cpu_to_fsm_m1_chipselect)))) & ((~pb_cpu_to_fsm_m1_qualified_request_ext_flash_1_s1 | ~(pb_cpu_to_fsm_m1_write & pb_cpu_to_fsm_m1_chipselect) | (1 & ((ext_flash_1_s1_wait_counter_eq_0 & ~d1_tb_fsm_avalon_slave_end_xfer)) & (pb_cpu_to_fsm_m1_dbs_address[1]) & (pb_cpu_to_fsm_m1_write & pb_cpu_to_fsm_m1_chipselect)))) & ((~pb_cpu_to_fsm_m1_qualified_request_ext_flash_s1 | ~(pb_cpu_to_fsm_m1_read & pb_cpu_to_fsm_m1_chipselect) | (1 & ((ext_flash_s1_wait_counter_eq_0 & ~d1_tb_fsm_avalon_slave_end_xfer)) & (pb_cpu_to_fsm_m1_dbs_address[1]) & (pb_cpu_to_fsm_m1_read & pb_cpu_to_fsm_m1_chipselect)))) & ((~pb_cpu_to_fsm_m1_qualified_request_ext_flash_s1 | ~(pb_cpu_to_fsm_m1_write & pb_cpu_to_fsm_m1_chipselect) | (1 & ((ext_flash_s1_wait_counter_eq_0 & ~d1_tb_fsm_avalon_slave_end_xfer)) & (pb_cpu_to_fsm_m1_dbs_address[1]) & (pb_cpu_to_fsm_m1_write & pb_cpu_to_fsm_m1_chipselect))));

  //cascaded wait assignment, which is an e_assign
  assign pb_cpu_to_fsm_m1_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign pb_cpu_to_fsm_m1_address_to_slave = pb_cpu_to_fsm_m1_address[25 : 0];

  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = (((~0) & pb_cpu_to_fsm_m1_requests_ext_flash_1_s1 & (pb_cpu_to_fsm_m1_write & pb_cpu_to_fsm_m1_chipselect) & !pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1)) |
    (((~0) & pb_cpu_to_fsm_m1_requests_ext_flash_s1 & (pb_cpu_to_fsm_m1_write & pb_cpu_to_fsm_m1_chipselect) & !pb_cpu_to_fsm_m1_byteenable_ext_flash_s1)) |
    ((pb_cpu_to_fsm_m1_granted_ext_flash_1_s1 & (pb_cpu_to_fsm_m1_read & pb_cpu_to_fsm_m1_chipselect) & 1 & 1 & ({ext_flash_1_s1_wait_counter_eq_0 & ~d1_tb_fsm_avalon_slave_end_xfer}))) |
    ((pb_cpu_to_fsm_m1_granted_ext_flash_1_s1 & (pb_cpu_to_fsm_m1_write & pb_cpu_to_fsm_m1_chipselect) & 1 & 1 & ({ext_flash_1_s1_wait_counter_eq_0 & ~d1_tb_fsm_avalon_slave_end_xfer}))) |
    ((pb_cpu_to_fsm_m1_granted_ext_flash_s1 & (pb_cpu_to_fsm_m1_read & pb_cpu_to_fsm_m1_chipselect) & 1 & 1 & ({ext_flash_s1_wait_counter_eq_0 & ~d1_tb_fsm_avalon_slave_end_xfer}))) |
    ((pb_cpu_to_fsm_m1_granted_ext_flash_s1 & (pb_cpu_to_fsm_m1_write & pb_cpu_to_fsm_m1_chipselect) & 1 & 1 & ({ext_flash_s1_wait_counter_eq_0 & ~d1_tb_fsm_avalon_slave_end_xfer})));

  //pb_cpu_to_fsm_m1_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_m1_read_but_no_slave_selected <= 0;
      else 
        pb_cpu_to_fsm_m1_read_but_no_slave_selected <= (pb_cpu_to_fsm_m1_read & pb_cpu_to_fsm_m1_chipselect) & pb_cpu_to_fsm_m1_run & ~pb_cpu_to_fsm_m1_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign pb_cpu_to_fsm_m1_is_granted_some_slave = pb_cpu_to_fsm_m1_granted_ext_flash_1_s1 |
    pb_cpu_to_fsm_m1_granted_ext_flash_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_pb_cpu_to_fsm_m1_readdatavalid = (pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1 & dbs_rdv_counter_overflow) |
    (pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1 & dbs_rdv_counter_overflow);

  //latent slave read data valid which is not flushed, which is an e_mux
  assign pb_cpu_to_fsm_m1_readdatavalid = pb_cpu_to_fsm_m1_read_but_no_slave_selected |
    pre_flush_pb_cpu_to_fsm_m1_readdatavalid |
    pb_cpu_to_fsm_m1_read_but_no_slave_selected |
    pre_flush_pb_cpu_to_fsm_m1_readdatavalid;

  //input to latent dbs-16 stored 0, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_0 = (pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1)? incoming_tb_fsm_data_with_Xs_converted_to_0 :
    incoming_tb_fsm_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((pb_cpu_to_fsm_m1_dbs_rdv_counter[1]) == 0))
          dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
    end


  //pb_cpu_to_fsm/m1 readdata mux, which is an e_mux
  assign pb_cpu_to_fsm_m1_readdata = ({32 {~pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1}} | {incoming_tb_fsm_data_with_Xs_converted_to_0[15 : 0],
    dbs_latent_16_reg_segment_0}) &
    ({32 {~pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1}} | {incoming_tb_fsm_data_with_Xs_converted_to_0[15 : 0],
    dbs_latent_16_reg_segment_0});

  //mux write dbs 1, which is an e_mux
  assign pb_cpu_to_fsm_m1_dbs_write_16 = (pb_cpu_to_fsm_m1_dbs_address[1])? pb_cpu_to_fsm_m1_writedata[31 : 16] :
    (~(pb_cpu_to_fsm_m1_dbs_address[1]))? pb_cpu_to_fsm_m1_writedata[15 : 0] :
    (pb_cpu_to_fsm_m1_dbs_address[1])? pb_cpu_to_fsm_m1_writedata[31 : 16] :
    pb_cpu_to_fsm_m1_writedata[15 : 0];

  //actual waitrequest port, which is an e_assign
  assign pb_cpu_to_fsm_m1_waitrequest = ~pb_cpu_to_fsm_m1_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_m1_latency_counter <= 0;
      else 
        pb_cpu_to_fsm_m1_latency_counter <= p1_pb_cpu_to_fsm_m1_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_pb_cpu_to_fsm_m1_latency_counter = ((pb_cpu_to_fsm_m1_run & (pb_cpu_to_fsm_m1_read & pb_cpu_to_fsm_m1_chipselect)))? latency_load_value :
    (pb_cpu_to_fsm_m1_latency_counter)? pb_cpu_to_fsm_m1_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({2 {pb_cpu_to_fsm_m1_requests_ext_flash_1_s1}} & 2) |
    ({2 {pb_cpu_to_fsm_m1_requests_ext_flash_s1}} & 2);

  //dbs count increment, which is an e_mux
  assign pb_cpu_to_fsm_m1_dbs_increment = (pb_cpu_to_fsm_m1_requests_ext_flash_1_s1)? 2 :
    (pb_cpu_to_fsm_m1_requests_ext_flash_s1)? 2 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = pb_cpu_to_fsm_m1_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = pb_cpu_to_fsm_m1_dbs_address + pb_cpu_to_fsm_m1_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_m1_dbs_address <= 0;
      else if (dbs_count_enable)
          pb_cpu_to_fsm_m1_dbs_address <= next_dbs_address;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign pb_cpu_to_fsm_m1_next_dbs_rdv_counter = pb_cpu_to_fsm_m1_dbs_rdv_counter + pb_cpu_to_fsm_m1_dbs_rdv_counter_inc;

  //pb_cpu_to_fsm_m1_rdv_inc_mux, which is an e_mux
  assign pb_cpu_to_fsm_m1_dbs_rdv_counter_inc = (pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1)? 2 :
    2;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1 |
    pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_m1_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          pb_cpu_to_fsm_m1_dbs_rdv_counter <= pb_cpu_to_fsm_m1_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = pb_cpu_to_fsm_m1_dbs_rdv_counter[1] & ~pb_cpu_to_fsm_m1_next_dbs_rdv_counter[1];


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pb_cpu_to_fsm_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_m1_address_last_time <= 0;
      else 
        pb_cpu_to_fsm_m1_address_last_time <= pb_cpu_to_fsm_m1_address;
    end


  //pb_cpu_to_fsm/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= pb_cpu_to_fsm_m1_waitrequest & pb_cpu_to_fsm_m1_chipselect;
    end


  //pb_cpu_to_fsm_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_fsm_m1_address != pb_cpu_to_fsm_m1_address_last_time))
        begin
          $write("%0d ns: pb_cpu_to_fsm_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_fsm_m1_chipselect check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_m1_chipselect_last_time <= 0;
      else 
        pb_cpu_to_fsm_m1_chipselect_last_time <= pb_cpu_to_fsm_m1_chipselect;
    end


  //pb_cpu_to_fsm_m1_chipselect matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_fsm_m1_chipselect != pb_cpu_to_fsm_m1_chipselect_last_time))
        begin
          $write("%0d ns: pb_cpu_to_fsm_m1_chipselect did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_fsm_m1_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_m1_burstcount_last_time <= 0;
      else 
        pb_cpu_to_fsm_m1_burstcount_last_time <= pb_cpu_to_fsm_m1_burstcount;
    end


  //pb_cpu_to_fsm_m1_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_fsm_m1_burstcount != pb_cpu_to_fsm_m1_burstcount_last_time))
        begin
          $write("%0d ns: pb_cpu_to_fsm_m1_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_fsm_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_m1_byteenable_last_time <= 0;
      else 
        pb_cpu_to_fsm_m1_byteenable_last_time <= pb_cpu_to_fsm_m1_byteenable;
    end


  //pb_cpu_to_fsm_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_fsm_m1_byteenable != pb_cpu_to_fsm_m1_byteenable_last_time))
        begin
          $write("%0d ns: pb_cpu_to_fsm_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_fsm_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_m1_read_last_time <= 0;
      else 
        pb_cpu_to_fsm_m1_read_last_time <= pb_cpu_to_fsm_m1_read;
    end


  //pb_cpu_to_fsm_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_fsm_m1_read != pb_cpu_to_fsm_m1_read_last_time))
        begin
          $write("%0d ns: pb_cpu_to_fsm_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_fsm_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_m1_write_last_time <= 0;
      else 
        pb_cpu_to_fsm_m1_write_last_time <= pb_cpu_to_fsm_m1_write;
    end


  //pb_cpu_to_fsm_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_fsm_m1_write != pb_cpu_to_fsm_m1_write_last_time))
        begin
          $write("%0d ns: pb_cpu_to_fsm_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_fsm_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_m1_writedata_last_time <= 0;
      else 
        pb_cpu_to_fsm_m1_writedata_last_time <= pb_cpu_to_fsm_m1_writedata;
    end


  //pb_cpu_to_fsm_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_fsm_m1_writedata != pb_cpu_to_fsm_m1_writedata_last_time) & (pb_cpu_to_fsm_m1_write & pb_cpu_to_fsm_m1_chipselect))
        begin
          $write("%0d ns: pb_cpu_to_fsm_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pb_cpu_to_fsm_bridge_arbitrator 
;



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_pb_cpu_to_io_s1_module (
                                                                // inputs:
                                                                 clear_fifo,
                                                                 clk,
                                                                 data_in,
                                                                 read,
                                                                 reset_n,
                                                                 sync_reset,
                                                                 write,

                                                                // outputs:
                                                                 data_out,
                                                                 empty,
                                                                 fifo_contains_ones_n,
                                                                 full
                                                              )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  wire             full_3;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_2;
  assign empty = !full_0;
  assign full_3 = 0;
  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    0;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pb_cpu_to_io_s1_arbitrator (
                                    // inputs:
                                     clk,
                                     cpu_data_master_address_to_slave,
                                     cpu_data_master_byteenable,
                                     cpu_data_master_debugaccess,
                                     cpu_data_master_latency_counter,
                                     cpu_data_master_read,
                                     cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register,
                                     cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register,
                                     cpu_data_master_write,
                                     cpu_data_master_writedata,
                                     pb_cpu_to_io_s1_endofpacket,
                                     pb_cpu_to_io_s1_readdata,
                                     pb_cpu_to_io_s1_readdatavalid,
                                     pb_cpu_to_io_s1_waitrequest,
                                     reset_n,

                                    // outputs:
                                     cpu_data_master_granted_pb_cpu_to_io_s1,
                                     cpu_data_master_qualified_request_pb_cpu_to_io_s1,
                                     cpu_data_master_read_data_valid_pb_cpu_to_io_s1,
                                     cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register,
                                     cpu_data_master_requests_pb_cpu_to_io_s1,
                                     d1_pb_cpu_to_io_s1_end_xfer,
                                     pb_cpu_to_io_s1_address,
                                     pb_cpu_to_io_s1_arbiterlock,
                                     pb_cpu_to_io_s1_arbiterlock2,
                                     pb_cpu_to_io_s1_burstcount,
                                     pb_cpu_to_io_s1_byteenable,
                                     pb_cpu_to_io_s1_chipselect,
                                     pb_cpu_to_io_s1_debugaccess,
                                     pb_cpu_to_io_s1_endofpacket_from_sa,
                                     pb_cpu_to_io_s1_nativeaddress,
                                     pb_cpu_to_io_s1_read,
                                     pb_cpu_to_io_s1_readdata_from_sa,
                                     pb_cpu_to_io_s1_reset_n,
                                     pb_cpu_to_io_s1_waitrequest_from_sa,
                                     pb_cpu_to_io_s1_write,
                                     pb_cpu_to_io_s1_writedata
                                  )
;

  output           cpu_data_master_granted_pb_cpu_to_io_s1;
  output           cpu_data_master_qualified_request_pb_cpu_to_io_s1;
  output           cpu_data_master_read_data_valid_pb_cpu_to_io_s1;
  output           cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register;
  output           cpu_data_master_requests_pb_cpu_to_io_s1;
  output           d1_pb_cpu_to_io_s1_end_xfer;
  output  [ 20: 0] pb_cpu_to_io_s1_address;
  output           pb_cpu_to_io_s1_arbiterlock;
  output           pb_cpu_to_io_s1_arbiterlock2;
  output           pb_cpu_to_io_s1_burstcount;
  output  [  3: 0] pb_cpu_to_io_s1_byteenable;
  output           pb_cpu_to_io_s1_chipselect;
  output           pb_cpu_to_io_s1_debugaccess;
  output           pb_cpu_to_io_s1_endofpacket_from_sa;
  output  [ 20: 0] pb_cpu_to_io_s1_nativeaddress;
  output           pb_cpu_to_io_s1_read;
  output  [ 31: 0] pb_cpu_to_io_s1_readdata_from_sa;
  output           pb_cpu_to_io_s1_reset_n;
  output           pb_cpu_to_io_s1_waitrequest_from_sa;
  output           pb_cpu_to_io_s1_write;
  output  [ 31: 0] pb_cpu_to_io_s1_writedata;
  input            clk;
  input   [ 28: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register;
  input            cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            pb_cpu_to_io_s1_endofpacket;
  input   [ 31: 0] pb_cpu_to_io_s1_readdata;
  input            pb_cpu_to_io_s1_readdatavalid;
  input            pb_cpu_to_io_s1_waitrequest;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_pb_cpu_to_io_s1;
  wire             cpu_data_master_qualified_request_pb_cpu_to_io_s1;
  wire             cpu_data_master_rdv_fifo_empty_pb_cpu_to_io_s1;
  wire             cpu_data_master_rdv_fifo_output_from_pb_cpu_to_io_s1;
  wire             cpu_data_master_read_data_valid_pb_cpu_to_io_s1;
  wire             cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register;
  wire             cpu_data_master_requests_pb_cpu_to_io_s1;
  wire             cpu_data_master_saved_grant_pb_cpu_to_io_s1;
  reg              d1_pb_cpu_to_io_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_pb_cpu_to_io_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 20: 0] pb_cpu_to_io_s1_address;
  wire             pb_cpu_to_io_s1_allgrants;
  wire             pb_cpu_to_io_s1_allow_new_arb_cycle;
  wire             pb_cpu_to_io_s1_any_bursting_master_saved_grant;
  wire             pb_cpu_to_io_s1_any_continuerequest;
  wire             pb_cpu_to_io_s1_arb_counter_enable;
  reg              pb_cpu_to_io_s1_arb_share_counter;
  wire             pb_cpu_to_io_s1_arb_share_counter_next_value;
  wire             pb_cpu_to_io_s1_arb_share_set_values;
  wire             pb_cpu_to_io_s1_arbiterlock;
  wire             pb_cpu_to_io_s1_arbiterlock2;
  wire             pb_cpu_to_io_s1_arbitration_holdoff_internal;
  wire             pb_cpu_to_io_s1_beginbursttransfer_internal;
  wire             pb_cpu_to_io_s1_begins_xfer;
  wire             pb_cpu_to_io_s1_burstcount;
  wire    [  3: 0] pb_cpu_to_io_s1_byteenable;
  wire             pb_cpu_to_io_s1_chipselect;
  wire             pb_cpu_to_io_s1_debugaccess;
  wire             pb_cpu_to_io_s1_end_xfer;
  wire             pb_cpu_to_io_s1_endofpacket_from_sa;
  wire             pb_cpu_to_io_s1_firsttransfer;
  wire             pb_cpu_to_io_s1_grant_vector;
  wire             pb_cpu_to_io_s1_in_a_read_cycle;
  wire             pb_cpu_to_io_s1_in_a_write_cycle;
  wire             pb_cpu_to_io_s1_master_qreq_vector;
  wire             pb_cpu_to_io_s1_move_on_to_next_transaction;
  wire    [ 20: 0] pb_cpu_to_io_s1_nativeaddress;
  wire             pb_cpu_to_io_s1_non_bursting_master_requests;
  wire             pb_cpu_to_io_s1_read;
  wire    [ 31: 0] pb_cpu_to_io_s1_readdata_from_sa;
  wire             pb_cpu_to_io_s1_readdatavalid_from_sa;
  reg              pb_cpu_to_io_s1_reg_firsttransfer;
  wire             pb_cpu_to_io_s1_reset_n;
  reg              pb_cpu_to_io_s1_slavearbiterlockenable;
  wire             pb_cpu_to_io_s1_slavearbiterlockenable2;
  wire             pb_cpu_to_io_s1_unreg_firsttransfer;
  wire             pb_cpu_to_io_s1_waitrequest_from_sa;
  wire             pb_cpu_to_io_s1_waits_for_read;
  wire             pb_cpu_to_io_s1_waits_for_write;
  wire             pb_cpu_to_io_s1_write;
  wire    [ 31: 0] pb_cpu_to_io_s1_writedata;
  wire    [ 28: 0] shifted_address_to_pb_cpu_to_io_s1_from_cpu_data_master;
  wire             wait_for_pb_cpu_to_io_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~pb_cpu_to_io_s1_end_xfer;
    end


  assign pb_cpu_to_io_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_pb_cpu_to_io_s1));
  //assign pb_cpu_to_io_s1_readdatavalid_from_sa = pb_cpu_to_io_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_cpu_to_io_s1_readdatavalid_from_sa = pb_cpu_to_io_s1_readdatavalid;

  //assign pb_cpu_to_io_s1_readdata_from_sa = pb_cpu_to_io_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_cpu_to_io_s1_readdata_from_sa = pb_cpu_to_io_s1_readdata;

  assign cpu_data_master_requests_pb_cpu_to_io_s1 = ({cpu_data_master_address_to_slave[28 : 23] , 23'b0} == 29'h8000000) & (cpu_data_master_read | cpu_data_master_write);
  //assign pb_cpu_to_io_s1_waitrequest_from_sa = pb_cpu_to_io_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_cpu_to_io_s1_waitrequest_from_sa = pb_cpu_to_io_s1_waitrequest;

  //pb_cpu_to_io_s1_arb_share_counter set values, which is an e_mux
  assign pb_cpu_to_io_s1_arb_share_set_values = 1;

  //pb_cpu_to_io_s1_non_bursting_master_requests mux, which is an e_mux
  assign pb_cpu_to_io_s1_non_bursting_master_requests = cpu_data_master_requests_pb_cpu_to_io_s1 |
    cpu_data_master_requests_pb_cpu_to_io_s1;

  //pb_cpu_to_io_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign pb_cpu_to_io_s1_any_bursting_master_saved_grant = 0;

  //pb_cpu_to_io_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign pb_cpu_to_io_s1_arb_share_counter_next_value = pb_cpu_to_io_s1_firsttransfer ? (pb_cpu_to_io_s1_arb_share_set_values - 1) : |pb_cpu_to_io_s1_arb_share_counter ? (pb_cpu_to_io_s1_arb_share_counter - 1) : 0;

  //pb_cpu_to_io_s1_allgrants all slave grants, which is an e_mux
  assign pb_cpu_to_io_s1_allgrants = (|pb_cpu_to_io_s1_grant_vector) |
    (|pb_cpu_to_io_s1_grant_vector);

  //pb_cpu_to_io_s1_end_xfer assignment, which is an e_assign
  assign pb_cpu_to_io_s1_end_xfer = ~(pb_cpu_to_io_s1_waits_for_read | pb_cpu_to_io_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_pb_cpu_to_io_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_pb_cpu_to_io_s1 = pb_cpu_to_io_s1_end_xfer & (~pb_cpu_to_io_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //pb_cpu_to_io_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign pb_cpu_to_io_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_pb_cpu_to_io_s1 & pb_cpu_to_io_s1_allgrants) | (end_xfer_arb_share_counter_term_pb_cpu_to_io_s1 & ~pb_cpu_to_io_s1_non_bursting_master_requests);

  //pb_cpu_to_io_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_io_s1_arb_share_counter <= 0;
      else if (pb_cpu_to_io_s1_arb_counter_enable)
          pb_cpu_to_io_s1_arb_share_counter <= pb_cpu_to_io_s1_arb_share_counter_next_value;
    end


  //pb_cpu_to_io_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_io_s1_slavearbiterlockenable <= 0;
      else if ((|pb_cpu_to_io_s1_master_qreq_vector & end_xfer_arb_share_counter_term_pb_cpu_to_io_s1) | (end_xfer_arb_share_counter_term_pb_cpu_to_io_s1 & ~pb_cpu_to_io_s1_non_bursting_master_requests))
          pb_cpu_to_io_s1_slavearbiterlockenable <= |pb_cpu_to_io_s1_arb_share_counter_next_value;
    end


  //cpu/data_master pb_cpu_to_io/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = pb_cpu_to_io_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //pb_cpu_to_io_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign pb_cpu_to_io_s1_slavearbiterlockenable2 = |pb_cpu_to_io_s1_arb_share_counter_next_value;

  //cpu/data_master pb_cpu_to_io/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = pb_cpu_to_io_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //pb_cpu_to_io_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign pb_cpu_to_io_s1_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_pb_cpu_to_io_s1 = cpu_data_master_requests_pb_cpu_to_io_s1 & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register) | (|cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register))));
  //unique name for pb_cpu_to_io_s1_move_on_to_next_transaction, which is an e_assign
  assign pb_cpu_to_io_s1_move_on_to_next_transaction = pb_cpu_to_io_s1_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_pb_cpu_to_io_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_pb_cpu_to_io_s1_module rdv_fifo_for_cpu_data_master_to_pb_cpu_to_io_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_pb_cpu_to_io_s1),
      .data_out             (cpu_data_master_rdv_fifo_output_from_pb_cpu_to_io_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_pb_cpu_to_io_s1),
      .full                 (),
      .read                 (pb_cpu_to_io_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~pb_cpu_to_io_s1_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register = ~cpu_data_master_rdv_fifo_empty_pb_cpu_to_io_s1;
  //local readdatavalid cpu_data_master_read_data_valid_pb_cpu_to_io_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_pb_cpu_to_io_s1 = pb_cpu_to_io_s1_readdatavalid_from_sa;

  //pb_cpu_to_io_s1_writedata mux, which is an e_mux
  assign pb_cpu_to_io_s1_writedata = cpu_data_master_writedata;

  //assign pb_cpu_to_io_s1_endofpacket_from_sa = pb_cpu_to_io_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_cpu_to_io_s1_endofpacket_from_sa = pb_cpu_to_io_s1_endofpacket;

  //master is always granted when requested
  assign cpu_data_master_granted_pb_cpu_to_io_s1 = cpu_data_master_qualified_request_pb_cpu_to_io_s1;

  //cpu/data_master saved-grant pb_cpu_to_io/s1, which is an e_assign
  assign cpu_data_master_saved_grant_pb_cpu_to_io_s1 = cpu_data_master_requests_pb_cpu_to_io_s1;

  //allow new arb cycle for pb_cpu_to_io/s1, which is an e_assign
  assign pb_cpu_to_io_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign pb_cpu_to_io_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign pb_cpu_to_io_s1_master_qreq_vector = 1;

  //pb_cpu_to_io_s1_reset_n assignment, which is an e_assign
  assign pb_cpu_to_io_s1_reset_n = reset_n;

  assign pb_cpu_to_io_s1_chipselect = cpu_data_master_granted_pb_cpu_to_io_s1;
  //pb_cpu_to_io_s1_firsttransfer first transaction, which is an e_assign
  assign pb_cpu_to_io_s1_firsttransfer = pb_cpu_to_io_s1_begins_xfer ? pb_cpu_to_io_s1_unreg_firsttransfer : pb_cpu_to_io_s1_reg_firsttransfer;

  //pb_cpu_to_io_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign pb_cpu_to_io_s1_unreg_firsttransfer = ~(pb_cpu_to_io_s1_slavearbiterlockenable & pb_cpu_to_io_s1_any_continuerequest);

  //pb_cpu_to_io_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_io_s1_reg_firsttransfer <= 1'b1;
      else if (pb_cpu_to_io_s1_begins_xfer)
          pb_cpu_to_io_s1_reg_firsttransfer <= pb_cpu_to_io_s1_unreg_firsttransfer;
    end


  //pb_cpu_to_io_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign pb_cpu_to_io_s1_beginbursttransfer_internal = pb_cpu_to_io_s1_begins_xfer;

  //pb_cpu_to_io_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign pb_cpu_to_io_s1_arbitration_holdoff_internal = pb_cpu_to_io_s1_begins_xfer & pb_cpu_to_io_s1_firsttransfer;

  //pb_cpu_to_io_s1_read assignment, which is an e_mux
  assign pb_cpu_to_io_s1_read = cpu_data_master_granted_pb_cpu_to_io_s1 & cpu_data_master_read;

  //pb_cpu_to_io_s1_write assignment, which is an e_mux
  assign pb_cpu_to_io_s1_write = cpu_data_master_granted_pb_cpu_to_io_s1 & cpu_data_master_write;

  assign shifted_address_to_pb_cpu_to_io_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //pb_cpu_to_io_s1_address mux, which is an e_mux
  assign pb_cpu_to_io_s1_address = shifted_address_to_pb_cpu_to_io_s1_from_cpu_data_master >> 2;

  //slaveid pb_cpu_to_io_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign pb_cpu_to_io_s1_nativeaddress = cpu_data_master_address_to_slave >> 2;

  //d1_pb_cpu_to_io_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_pb_cpu_to_io_s1_end_xfer <= 1;
      else 
        d1_pb_cpu_to_io_s1_end_xfer <= pb_cpu_to_io_s1_end_xfer;
    end


  //pb_cpu_to_io_s1_waits_for_read in a cycle, which is an e_mux
  assign pb_cpu_to_io_s1_waits_for_read = pb_cpu_to_io_s1_in_a_read_cycle & pb_cpu_to_io_s1_waitrequest_from_sa;

  //pb_cpu_to_io_s1_in_a_read_cycle assignment, which is an e_assign
  assign pb_cpu_to_io_s1_in_a_read_cycle = cpu_data_master_granted_pb_cpu_to_io_s1 & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = pb_cpu_to_io_s1_in_a_read_cycle;

  //pb_cpu_to_io_s1_waits_for_write in a cycle, which is an e_mux
  assign pb_cpu_to_io_s1_waits_for_write = pb_cpu_to_io_s1_in_a_write_cycle & pb_cpu_to_io_s1_waitrequest_from_sa;

  //pb_cpu_to_io_s1_in_a_write_cycle assignment, which is an e_assign
  assign pb_cpu_to_io_s1_in_a_write_cycle = cpu_data_master_granted_pb_cpu_to_io_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = pb_cpu_to_io_s1_in_a_write_cycle;

  assign wait_for_pb_cpu_to_io_s1_counter = 0;
  //pb_cpu_to_io_s1_byteenable byte enable port mux, which is an e_mux
  assign pb_cpu_to_io_s1_byteenable = (cpu_data_master_granted_pb_cpu_to_io_s1)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign pb_cpu_to_io_s1_burstcount = 1;

  //pb_cpu_to_io/s1 arbiterlock assigned from _handle_arbiterlock, which is an e_mux
  assign pb_cpu_to_io_s1_arbiterlock = cpu_data_master_arbiterlock;

  //pb_cpu_to_io/s1 arbiterlock2 assigned from _handle_arbiterlock2, which is an e_mux
  assign pb_cpu_to_io_s1_arbiterlock2 = cpu_data_master_arbiterlock2;

  //debugaccess mux, which is an e_mux
  assign pb_cpu_to_io_s1_debugaccess = (cpu_data_master_granted_pb_cpu_to_io_s1)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pb_cpu_to_io/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pb_cpu_to_io_m1_arbitrator (
                                    // inputs:
                                     button_pio_s1_readdata_from_sa,
                                     clk,
                                     d1_button_pio_s1_end_xfer,
                                     d1_descriptor_memory_s1_end_xfer,
                                     d1_dipsw_pio_s1_end_xfer,
                                     d1_jtag_uart_avalon_jtag_slave_end_xfer,
                                     d1_led_pio_s1_end_xfer,
                                     d1_sgdma_rx_csr_end_xfer,
                                     d1_sgdma_tx_csr_end_xfer,
                                     d1_sysid_control_slave_end_xfer,
                                     d1_timer_1ms_s1_end_xfer,
                                     d1_tse_mac_control_port_end_xfer,
                                     d1_uart_s1_end_xfer,
                                     descriptor_memory_s1_readdata_from_sa,
                                     dipsw_pio_s1_readdata_from_sa,
                                     jtag_uart_avalon_jtag_slave_readdata_from_sa,
                                     jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
                                     led_pio_s1_readdata_from_sa,
                                     pb_cpu_to_io_m1_address,
                                     pb_cpu_to_io_m1_burstcount,
                                     pb_cpu_to_io_m1_byteenable,
                                     pb_cpu_to_io_m1_chipselect,
                                     pb_cpu_to_io_m1_granted_button_pio_s1,
                                     pb_cpu_to_io_m1_granted_descriptor_memory_s1,
                                     pb_cpu_to_io_m1_granted_dipsw_pio_s1,
                                     pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave,
                                     pb_cpu_to_io_m1_granted_led_pio_s1,
                                     pb_cpu_to_io_m1_granted_sgdma_rx_csr,
                                     pb_cpu_to_io_m1_granted_sgdma_tx_csr,
                                     pb_cpu_to_io_m1_granted_sysid_control_slave,
                                     pb_cpu_to_io_m1_granted_timer_1ms_s1,
                                     pb_cpu_to_io_m1_granted_tse_mac_control_port,
                                     pb_cpu_to_io_m1_granted_uart_s1,
                                     pb_cpu_to_io_m1_qualified_request_button_pio_s1,
                                     pb_cpu_to_io_m1_qualified_request_descriptor_memory_s1,
                                     pb_cpu_to_io_m1_qualified_request_dipsw_pio_s1,
                                     pb_cpu_to_io_m1_qualified_request_jtag_uart_avalon_jtag_slave,
                                     pb_cpu_to_io_m1_qualified_request_led_pio_s1,
                                     pb_cpu_to_io_m1_qualified_request_sgdma_rx_csr,
                                     pb_cpu_to_io_m1_qualified_request_sgdma_tx_csr,
                                     pb_cpu_to_io_m1_qualified_request_sysid_control_slave,
                                     pb_cpu_to_io_m1_qualified_request_timer_1ms_s1,
                                     pb_cpu_to_io_m1_qualified_request_tse_mac_control_port,
                                     pb_cpu_to_io_m1_qualified_request_uart_s1,
                                     pb_cpu_to_io_m1_read,
                                     pb_cpu_to_io_m1_read_data_valid_button_pio_s1,
                                     pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1,
                                     pb_cpu_to_io_m1_read_data_valid_dipsw_pio_s1,
                                     pb_cpu_to_io_m1_read_data_valid_jtag_uart_avalon_jtag_slave,
                                     pb_cpu_to_io_m1_read_data_valid_led_pio_s1,
                                     pb_cpu_to_io_m1_read_data_valid_sgdma_rx_csr,
                                     pb_cpu_to_io_m1_read_data_valid_sgdma_tx_csr,
                                     pb_cpu_to_io_m1_read_data_valid_sysid_control_slave,
                                     pb_cpu_to_io_m1_read_data_valid_timer_1ms_s1,
                                     pb_cpu_to_io_m1_read_data_valid_tse_mac_control_port,
                                     pb_cpu_to_io_m1_read_data_valid_uart_s1,
                                     pb_cpu_to_io_m1_requests_button_pio_s1,
                                     pb_cpu_to_io_m1_requests_descriptor_memory_s1,
                                     pb_cpu_to_io_m1_requests_dipsw_pio_s1,
                                     pb_cpu_to_io_m1_requests_jtag_uart_avalon_jtag_slave,
                                     pb_cpu_to_io_m1_requests_led_pio_s1,
                                     pb_cpu_to_io_m1_requests_sgdma_rx_csr,
                                     pb_cpu_to_io_m1_requests_sgdma_tx_csr,
                                     pb_cpu_to_io_m1_requests_sysid_control_slave,
                                     pb_cpu_to_io_m1_requests_timer_1ms_s1,
                                     pb_cpu_to_io_m1_requests_tse_mac_control_port,
                                     pb_cpu_to_io_m1_requests_uart_s1,
                                     pb_cpu_to_io_m1_write,
                                     pb_cpu_to_io_m1_writedata,
                                     reset_n,
                                     sgdma_rx_csr_readdata_from_sa,
                                     sgdma_tx_csr_readdata_from_sa,
                                     sysid_control_slave_readdata_from_sa,
                                     timer_1ms_s1_readdata_from_sa,
                                     tse_mac_control_port_readdata_from_sa,
                                     tse_mac_control_port_waitrequest_from_sa,
                                     uart_s1_readdata_from_sa,

                                    // outputs:
                                     pb_cpu_to_io_m1_address_to_slave,
                                     pb_cpu_to_io_m1_latency_counter,
                                     pb_cpu_to_io_m1_readdata,
                                     pb_cpu_to_io_m1_readdatavalid,
                                     pb_cpu_to_io_m1_waitrequest
                                  )
;

  output  [ 22: 0] pb_cpu_to_io_m1_address_to_slave;
  output           pb_cpu_to_io_m1_latency_counter;
  output  [ 31: 0] pb_cpu_to_io_m1_readdata;
  output           pb_cpu_to_io_m1_readdatavalid;
  output           pb_cpu_to_io_m1_waitrequest;
  input   [  2: 0] button_pio_s1_readdata_from_sa;
  input            clk;
  input            d1_button_pio_s1_end_xfer;
  input            d1_descriptor_memory_s1_end_xfer;
  input            d1_dipsw_pio_s1_end_xfer;
  input            d1_jtag_uart_avalon_jtag_slave_end_xfer;
  input            d1_led_pio_s1_end_xfer;
  input            d1_sgdma_rx_csr_end_xfer;
  input            d1_sgdma_tx_csr_end_xfer;
  input            d1_sysid_control_slave_end_xfer;
  input            d1_timer_1ms_s1_end_xfer;
  input            d1_tse_mac_control_port_end_xfer;
  input            d1_uart_s1_end_xfer;
  input   [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  input   [  7: 0] dipsw_pio_s1_readdata_from_sa;
  input   [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  input            jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  input   [ 15: 0] led_pio_s1_readdata_from_sa;
  input   [ 22: 0] pb_cpu_to_io_m1_address;
  input            pb_cpu_to_io_m1_burstcount;
  input   [  3: 0] pb_cpu_to_io_m1_byteenable;
  input            pb_cpu_to_io_m1_chipselect;
  input            pb_cpu_to_io_m1_granted_button_pio_s1;
  input            pb_cpu_to_io_m1_granted_descriptor_memory_s1;
  input            pb_cpu_to_io_m1_granted_dipsw_pio_s1;
  input            pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave;
  input            pb_cpu_to_io_m1_granted_led_pio_s1;
  input            pb_cpu_to_io_m1_granted_sgdma_rx_csr;
  input            pb_cpu_to_io_m1_granted_sgdma_tx_csr;
  input            pb_cpu_to_io_m1_granted_sysid_control_slave;
  input            pb_cpu_to_io_m1_granted_timer_1ms_s1;
  input            pb_cpu_to_io_m1_granted_tse_mac_control_port;
  input            pb_cpu_to_io_m1_granted_uart_s1;
  input            pb_cpu_to_io_m1_qualified_request_button_pio_s1;
  input            pb_cpu_to_io_m1_qualified_request_descriptor_memory_s1;
  input            pb_cpu_to_io_m1_qualified_request_dipsw_pio_s1;
  input            pb_cpu_to_io_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  input            pb_cpu_to_io_m1_qualified_request_led_pio_s1;
  input            pb_cpu_to_io_m1_qualified_request_sgdma_rx_csr;
  input            pb_cpu_to_io_m1_qualified_request_sgdma_tx_csr;
  input            pb_cpu_to_io_m1_qualified_request_sysid_control_slave;
  input            pb_cpu_to_io_m1_qualified_request_timer_1ms_s1;
  input            pb_cpu_to_io_m1_qualified_request_tse_mac_control_port;
  input            pb_cpu_to_io_m1_qualified_request_uart_s1;
  input            pb_cpu_to_io_m1_read;
  input            pb_cpu_to_io_m1_read_data_valid_button_pio_s1;
  input            pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1;
  input            pb_cpu_to_io_m1_read_data_valid_dipsw_pio_s1;
  input            pb_cpu_to_io_m1_read_data_valid_jtag_uart_avalon_jtag_slave;
  input            pb_cpu_to_io_m1_read_data_valid_led_pio_s1;
  input            pb_cpu_to_io_m1_read_data_valid_sgdma_rx_csr;
  input            pb_cpu_to_io_m1_read_data_valid_sgdma_tx_csr;
  input            pb_cpu_to_io_m1_read_data_valid_sysid_control_slave;
  input            pb_cpu_to_io_m1_read_data_valid_timer_1ms_s1;
  input            pb_cpu_to_io_m1_read_data_valid_tse_mac_control_port;
  input            pb_cpu_to_io_m1_read_data_valid_uart_s1;
  input            pb_cpu_to_io_m1_requests_button_pio_s1;
  input            pb_cpu_to_io_m1_requests_descriptor_memory_s1;
  input            pb_cpu_to_io_m1_requests_dipsw_pio_s1;
  input            pb_cpu_to_io_m1_requests_jtag_uart_avalon_jtag_slave;
  input            pb_cpu_to_io_m1_requests_led_pio_s1;
  input            pb_cpu_to_io_m1_requests_sgdma_rx_csr;
  input            pb_cpu_to_io_m1_requests_sgdma_tx_csr;
  input            pb_cpu_to_io_m1_requests_sysid_control_slave;
  input            pb_cpu_to_io_m1_requests_timer_1ms_s1;
  input            pb_cpu_to_io_m1_requests_tse_mac_control_port;
  input            pb_cpu_to_io_m1_requests_uart_s1;
  input            pb_cpu_to_io_m1_write;
  input   [ 31: 0] pb_cpu_to_io_m1_writedata;
  input            reset_n;
  input   [ 31: 0] sgdma_rx_csr_readdata_from_sa;
  input   [ 31: 0] sgdma_tx_csr_readdata_from_sa;
  input   [ 31: 0] sysid_control_slave_readdata_from_sa;
  input   [ 15: 0] timer_1ms_s1_readdata_from_sa;
  input   [ 31: 0] tse_mac_control_port_readdata_from_sa;
  input            tse_mac_control_port_waitrequest_from_sa;
  input   [ 15: 0] uart_s1_readdata_from_sa;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_pb_cpu_to_io_m1_latency_counter;
  reg     [ 22: 0] pb_cpu_to_io_m1_address_last_time;
  wire    [ 22: 0] pb_cpu_to_io_m1_address_to_slave;
  reg              pb_cpu_to_io_m1_burstcount_last_time;
  reg     [  3: 0] pb_cpu_to_io_m1_byteenable_last_time;
  reg              pb_cpu_to_io_m1_chipselect_last_time;
  wire             pb_cpu_to_io_m1_is_granted_some_slave;
  reg              pb_cpu_to_io_m1_latency_counter;
  reg              pb_cpu_to_io_m1_read_but_no_slave_selected;
  reg              pb_cpu_to_io_m1_read_last_time;
  wire    [ 31: 0] pb_cpu_to_io_m1_readdata;
  wire             pb_cpu_to_io_m1_readdatavalid;
  wire             pb_cpu_to_io_m1_run;
  wire             pb_cpu_to_io_m1_waitrequest;
  reg              pb_cpu_to_io_m1_write_last_time;
  reg     [ 31: 0] pb_cpu_to_io_m1_writedata_last_time;
  wire             pre_flush_pb_cpu_to_io_m1_readdatavalid;
  wire             r_0;
  wire             r_1;
  wire             r_2;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (pb_cpu_to_io_m1_qualified_request_button_pio_s1 | ~pb_cpu_to_io_m1_requests_button_pio_s1) & ((~pb_cpu_to_io_m1_qualified_request_button_pio_s1 | ~(pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) | (1 & ~d1_button_pio_s1_end_xfer & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)))) & ((~pb_cpu_to_io_m1_qualified_request_button_pio_s1 | ~(pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect) | (1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect)))) & 1 & (pb_cpu_to_io_m1_qualified_request_descriptor_memory_s1 | ~pb_cpu_to_io_m1_requests_descriptor_memory_s1) & (pb_cpu_to_io_m1_granted_descriptor_memory_s1 | ~pb_cpu_to_io_m1_qualified_request_descriptor_memory_s1) & ((~pb_cpu_to_io_m1_qualified_request_descriptor_memory_s1 | ~pb_cpu_to_io_m1_chipselect | (1 & pb_cpu_to_io_m1_chipselect))) & ((~pb_cpu_to_io_m1_qualified_request_descriptor_memory_s1 | ~pb_cpu_to_io_m1_chipselect | (1 & pb_cpu_to_io_m1_chipselect))) & 1 & (pb_cpu_to_io_m1_qualified_request_dipsw_pio_s1 | ~pb_cpu_to_io_m1_requests_dipsw_pio_s1) & ((~pb_cpu_to_io_m1_qualified_request_dipsw_pio_s1 | ~(pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) | (1 & ~d1_dipsw_pio_s1_end_xfer & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)))) & ((~pb_cpu_to_io_m1_qualified_request_dipsw_pio_s1 | ~(pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect) | (1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect)))) & 1 & (pb_cpu_to_io_m1_qualified_request_jtag_uart_avalon_jtag_slave | ~pb_cpu_to_io_m1_requests_jtag_uart_avalon_jtag_slave) & ((~pb_cpu_to_io_m1_qualified_request_jtag_uart_avalon_jtag_slave | ~pb_cpu_to_io_m1_chipselect | (1 & ~jtag_uart_avalon_jtag_slave_waitrequest_from_sa & pb_cpu_to_io_m1_chipselect))) & ((~pb_cpu_to_io_m1_qualified_request_jtag_uart_avalon_jtag_slave | ~pb_cpu_to_io_m1_chipselect | (1 & ~jtag_uart_avalon_jtag_slave_waitrequest_from_sa & pb_cpu_to_io_m1_chipselect))) & 1 & (pb_cpu_to_io_m1_qualified_request_led_pio_s1 | ~pb_cpu_to_io_m1_requests_led_pio_s1) & ((~pb_cpu_to_io_m1_qualified_request_led_pio_s1 | ~(pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) | (1 & ~d1_led_pio_s1_end_xfer & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect))));

  //cascaded wait assignment, which is an e_assign
  assign pb_cpu_to_io_m1_run = r_0 & r_1 & r_2;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = ((~pb_cpu_to_io_m1_qualified_request_led_pio_s1 | ~(pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect) | (1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect)))) & 1 & (pb_cpu_to_io_m1_qualified_request_sgdma_rx_csr | ~pb_cpu_to_io_m1_requests_sgdma_rx_csr) & ((~pb_cpu_to_io_m1_qualified_request_sgdma_rx_csr | ~(pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) | (1 & ~d1_sgdma_rx_csr_end_xfer & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)))) & ((~pb_cpu_to_io_m1_qualified_request_sgdma_rx_csr | ~(pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect) | (1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect)))) & 1 & (pb_cpu_to_io_m1_qualified_request_sgdma_tx_csr | ~pb_cpu_to_io_m1_requests_sgdma_tx_csr) & ((~pb_cpu_to_io_m1_qualified_request_sgdma_tx_csr | ~(pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) | (1 & ~d1_sgdma_tx_csr_end_xfer & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)))) & ((~pb_cpu_to_io_m1_qualified_request_sgdma_tx_csr | ~(pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect) | (1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect)))) & 1 & (pb_cpu_to_io_m1_qualified_request_sysid_control_slave | ~pb_cpu_to_io_m1_requests_sysid_control_slave) & ((~pb_cpu_to_io_m1_qualified_request_sysid_control_slave | ~(pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) | (1 & ~d1_sysid_control_slave_end_xfer & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)))) & ((~pb_cpu_to_io_m1_qualified_request_sysid_control_slave | ~(pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect) | (1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect)))) & 1 & (pb_cpu_to_io_m1_qualified_request_timer_1ms_s1 | ~pb_cpu_to_io_m1_requests_timer_1ms_s1) & ((~pb_cpu_to_io_m1_qualified_request_timer_1ms_s1 | ~(pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) | (1 & ~d1_timer_1ms_s1_end_xfer & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)))) & ((~pb_cpu_to_io_m1_qualified_request_timer_1ms_s1 | ~(pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect) | (1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect)))) & 1 & (pb_cpu_to_io_m1_qualified_request_tse_mac_control_port | ~pb_cpu_to_io_m1_requests_tse_mac_control_port) & ((~pb_cpu_to_io_m1_qualified_request_tse_mac_control_port | ~pb_cpu_to_io_m1_chipselect | (1 & ~tse_mac_control_port_waitrequest_from_sa & pb_cpu_to_io_m1_chipselect)));

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = ((~pb_cpu_to_io_m1_qualified_request_tse_mac_control_port | ~pb_cpu_to_io_m1_chipselect | (1 & ~tse_mac_control_port_waitrequest_from_sa & pb_cpu_to_io_m1_chipselect))) & 1 & (pb_cpu_to_io_m1_qualified_request_uart_s1 | ~pb_cpu_to_io_m1_requests_uart_s1) & ((~pb_cpu_to_io_m1_qualified_request_uart_s1 | ~pb_cpu_to_io_m1_chipselect | (1 & ~d1_uart_s1_end_xfer & pb_cpu_to_io_m1_chipselect))) & ((~pb_cpu_to_io_m1_qualified_request_uart_s1 | ~pb_cpu_to_io_m1_chipselect | (1 & ~d1_uart_s1_end_xfer & pb_cpu_to_io_m1_chipselect)));

  //optimize select-logic by passing only those address bits which matter.
  assign pb_cpu_to_io_m1_address_to_slave = {pb_cpu_to_io_m1_address[22],
    7'b0,
    pb_cpu_to_io_m1_address[14 : 0]};

  //pb_cpu_to_io_m1_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_io_m1_read_but_no_slave_selected <= 0;
      else 
        pb_cpu_to_io_m1_read_but_no_slave_selected <= (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & pb_cpu_to_io_m1_run & ~pb_cpu_to_io_m1_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign pb_cpu_to_io_m1_is_granted_some_slave = pb_cpu_to_io_m1_granted_button_pio_s1 |
    pb_cpu_to_io_m1_granted_descriptor_memory_s1 |
    pb_cpu_to_io_m1_granted_dipsw_pio_s1 |
    pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave |
    pb_cpu_to_io_m1_granted_led_pio_s1 |
    pb_cpu_to_io_m1_granted_sgdma_rx_csr |
    pb_cpu_to_io_m1_granted_sgdma_tx_csr |
    pb_cpu_to_io_m1_granted_sysid_control_slave |
    pb_cpu_to_io_m1_granted_timer_1ms_s1 |
    pb_cpu_to_io_m1_granted_tse_mac_control_port |
    pb_cpu_to_io_m1_granted_uart_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_pb_cpu_to_io_m1_readdatavalid = pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign pb_cpu_to_io_m1_readdatavalid = pb_cpu_to_io_m1_read_but_no_slave_selected |
    pre_flush_pb_cpu_to_io_m1_readdatavalid |
    pb_cpu_to_io_m1_read_data_valid_button_pio_s1 |
    pb_cpu_to_io_m1_read_but_no_slave_selected |
    pre_flush_pb_cpu_to_io_m1_readdatavalid |
    pb_cpu_to_io_m1_read_but_no_slave_selected |
    pre_flush_pb_cpu_to_io_m1_readdatavalid |
    pb_cpu_to_io_m1_read_data_valid_dipsw_pio_s1 |
    pb_cpu_to_io_m1_read_but_no_slave_selected |
    pre_flush_pb_cpu_to_io_m1_readdatavalid |
    pb_cpu_to_io_m1_read_data_valid_jtag_uart_avalon_jtag_slave |
    pb_cpu_to_io_m1_read_but_no_slave_selected |
    pre_flush_pb_cpu_to_io_m1_readdatavalid |
    pb_cpu_to_io_m1_read_data_valid_led_pio_s1 |
    pb_cpu_to_io_m1_read_but_no_slave_selected |
    pre_flush_pb_cpu_to_io_m1_readdatavalid |
    pb_cpu_to_io_m1_read_data_valid_sgdma_rx_csr |
    pb_cpu_to_io_m1_read_but_no_slave_selected |
    pre_flush_pb_cpu_to_io_m1_readdatavalid |
    pb_cpu_to_io_m1_read_data_valid_sgdma_tx_csr |
    pb_cpu_to_io_m1_read_but_no_slave_selected |
    pre_flush_pb_cpu_to_io_m1_readdatavalid |
    pb_cpu_to_io_m1_read_data_valid_sysid_control_slave |
    pb_cpu_to_io_m1_read_but_no_slave_selected |
    pre_flush_pb_cpu_to_io_m1_readdatavalid |
    pb_cpu_to_io_m1_read_data_valid_timer_1ms_s1 |
    pb_cpu_to_io_m1_read_but_no_slave_selected |
    pre_flush_pb_cpu_to_io_m1_readdatavalid |
    pb_cpu_to_io_m1_read_data_valid_tse_mac_control_port |
    pb_cpu_to_io_m1_read_but_no_slave_selected |
    pre_flush_pb_cpu_to_io_m1_readdatavalid |
    pb_cpu_to_io_m1_read_data_valid_uart_s1;

  //pb_cpu_to_io/m1 readdata mux, which is an e_mux
  assign pb_cpu_to_io_m1_readdata = ({32 {~((pb_cpu_to_io_m1_qualified_request_button_pio_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)))}} | button_pio_s1_readdata_from_sa) &
    ({32 {~pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1}} | descriptor_memory_s1_readdata_from_sa) &
    ({32 {~((pb_cpu_to_io_m1_qualified_request_dipsw_pio_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)))}} | dipsw_pio_s1_readdata_from_sa) &
    ({32 {~((pb_cpu_to_io_m1_qualified_request_jtag_uart_avalon_jtag_slave & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)))}} | jtag_uart_avalon_jtag_slave_readdata_from_sa) &
    ({32 {~((pb_cpu_to_io_m1_qualified_request_led_pio_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)))}} | led_pio_s1_readdata_from_sa) &
    ({32 {~((pb_cpu_to_io_m1_qualified_request_sgdma_rx_csr & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)))}} | sgdma_rx_csr_readdata_from_sa) &
    ({32 {~((pb_cpu_to_io_m1_qualified_request_sgdma_tx_csr & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)))}} | sgdma_tx_csr_readdata_from_sa) &
    ({32 {~((pb_cpu_to_io_m1_qualified_request_sysid_control_slave & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)))}} | sysid_control_slave_readdata_from_sa) &
    ({32 {~((pb_cpu_to_io_m1_qualified_request_timer_1ms_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)))}} | timer_1ms_s1_readdata_from_sa) &
    ({32 {~((pb_cpu_to_io_m1_qualified_request_tse_mac_control_port & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)))}} | tse_mac_control_port_readdata_from_sa) &
    ({32 {~((pb_cpu_to_io_m1_qualified_request_uart_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)))}} | uart_s1_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign pb_cpu_to_io_m1_waitrequest = ~pb_cpu_to_io_m1_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_io_m1_latency_counter <= 0;
      else 
        pb_cpu_to_io_m1_latency_counter <= p1_pb_cpu_to_io_m1_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_pb_cpu_to_io_m1_latency_counter = ((pb_cpu_to_io_m1_run & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect)))? latency_load_value :
    (pb_cpu_to_io_m1_latency_counter)? pb_cpu_to_io_m1_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {1 {pb_cpu_to_io_m1_requests_descriptor_memory_s1}} & 1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pb_cpu_to_io_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_io_m1_address_last_time <= 0;
      else 
        pb_cpu_to_io_m1_address_last_time <= pb_cpu_to_io_m1_address;
    end


  //pb_cpu_to_io/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= pb_cpu_to_io_m1_waitrequest & pb_cpu_to_io_m1_chipselect;
    end


  //pb_cpu_to_io_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_io_m1_address != pb_cpu_to_io_m1_address_last_time))
        begin
          $write("%0d ns: pb_cpu_to_io_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_io_m1_chipselect check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_io_m1_chipselect_last_time <= 0;
      else 
        pb_cpu_to_io_m1_chipselect_last_time <= pb_cpu_to_io_m1_chipselect;
    end


  //pb_cpu_to_io_m1_chipselect matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_io_m1_chipselect != pb_cpu_to_io_m1_chipselect_last_time))
        begin
          $write("%0d ns: pb_cpu_to_io_m1_chipselect did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_io_m1_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_io_m1_burstcount_last_time <= 0;
      else 
        pb_cpu_to_io_m1_burstcount_last_time <= pb_cpu_to_io_m1_burstcount;
    end


  //pb_cpu_to_io_m1_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_io_m1_burstcount != pb_cpu_to_io_m1_burstcount_last_time))
        begin
          $write("%0d ns: pb_cpu_to_io_m1_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_io_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_io_m1_byteenable_last_time <= 0;
      else 
        pb_cpu_to_io_m1_byteenable_last_time <= pb_cpu_to_io_m1_byteenable;
    end


  //pb_cpu_to_io_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_io_m1_byteenable != pb_cpu_to_io_m1_byteenable_last_time))
        begin
          $write("%0d ns: pb_cpu_to_io_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_io_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_io_m1_read_last_time <= 0;
      else 
        pb_cpu_to_io_m1_read_last_time <= pb_cpu_to_io_m1_read;
    end


  //pb_cpu_to_io_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_io_m1_read != pb_cpu_to_io_m1_read_last_time))
        begin
          $write("%0d ns: pb_cpu_to_io_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_io_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_io_m1_write_last_time <= 0;
      else 
        pb_cpu_to_io_m1_write_last_time <= pb_cpu_to_io_m1_write;
    end


  //pb_cpu_to_io_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_io_m1_write != pb_cpu_to_io_m1_write_last_time))
        begin
          $write("%0d ns: pb_cpu_to_io_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_cpu_to_io_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_io_m1_writedata_last_time <= 0;
      else 
        pb_cpu_to_io_m1_writedata_last_time <= pb_cpu_to_io_m1_writedata;
    end


  //pb_cpu_to_io_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_cpu_to_io_m1_writedata != pb_cpu_to_io_m1_writedata_last_time) & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect))
        begin
          $write("%0d ns: pb_cpu_to_io_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pb_cpu_to_io_bridge_arbitrator 
;



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_sgdma_tx_m_read_to_pb_dma_to_ddr3_top_s1_module (
                                                                      // inputs:
                                                                       clear_fifo,
                                                                       clk,
                                                                       data_in,
                                                                       read,
                                                                       reset_n,
                                                                       sync_reset,
                                                                       write,

                                                                      // outputs:
                                                                       data_out,
                                                                       empty,
                                                                       fifo_contains_ones_n,
                                                                       full
                                                                    )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  wire             full_34;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_33;
  assign empty = !full_0;
  assign full_34 = 0;
  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    0;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pb_dma_to_ddr3_top_s1_arbitrator (
                                          // inputs:
                                           clk,
                                           pb_dma_to_ddr3_top_s1_endofpacket,
                                           pb_dma_to_ddr3_top_s1_readdata,
                                           pb_dma_to_ddr3_top_s1_readdatavalid,
                                           pb_dma_to_ddr3_top_s1_waitrequest,
                                           reset_n,
                                           sgdma_rx_m_write_address_to_slave,
                                           sgdma_rx_m_write_byteenable,
                                           sgdma_rx_m_write_write,
                                           sgdma_rx_m_write_writedata,
                                           sgdma_tx_m_read_address_to_slave,
                                           sgdma_tx_m_read_latency_counter,
                                           sgdma_tx_m_read_read,

                                          // outputs:
                                           d1_pb_dma_to_ddr3_top_s1_end_xfer,
                                           pb_dma_to_ddr3_top_s1_address,
                                           pb_dma_to_ddr3_top_s1_arbiterlock,
                                           pb_dma_to_ddr3_top_s1_arbiterlock2,
                                           pb_dma_to_ddr3_top_s1_burstcount,
                                           pb_dma_to_ddr3_top_s1_byteenable,
                                           pb_dma_to_ddr3_top_s1_chipselect,
                                           pb_dma_to_ddr3_top_s1_debugaccess,
                                           pb_dma_to_ddr3_top_s1_endofpacket_from_sa,
                                           pb_dma_to_ddr3_top_s1_nativeaddress,
                                           pb_dma_to_ddr3_top_s1_read,
                                           pb_dma_to_ddr3_top_s1_readdata_from_sa,
                                           pb_dma_to_ddr3_top_s1_reset_n,
                                           pb_dma_to_ddr3_top_s1_waitrequest_from_sa,
                                           pb_dma_to_ddr3_top_s1_write,
                                           pb_dma_to_ddr3_top_s1_writedata,
                                           sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1,
                                           sgdma_rx_m_write_qualified_request_pb_dma_to_ddr3_top_s1,
                                           sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1,
                                           sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1,
                                           sgdma_tx_m_read_qualified_request_pb_dma_to_ddr3_top_s1,
                                           sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1,
                                           sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1_shift_register,
                                           sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1
                                        )
;

  output           d1_pb_dma_to_ddr3_top_s1_end_xfer;
  output  [ 24: 0] pb_dma_to_ddr3_top_s1_address;
  output           pb_dma_to_ddr3_top_s1_arbiterlock;
  output           pb_dma_to_ddr3_top_s1_arbiterlock2;
  output           pb_dma_to_ddr3_top_s1_burstcount;
  output  [  3: 0] pb_dma_to_ddr3_top_s1_byteenable;
  output           pb_dma_to_ddr3_top_s1_chipselect;
  output           pb_dma_to_ddr3_top_s1_debugaccess;
  output           pb_dma_to_ddr3_top_s1_endofpacket_from_sa;
  output  [ 24: 0] pb_dma_to_ddr3_top_s1_nativeaddress;
  output           pb_dma_to_ddr3_top_s1_read;
  output  [ 31: 0] pb_dma_to_ddr3_top_s1_readdata_from_sa;
  output           pb_dma_to_ddr3_top_s1_reset_n;
  output           pb_dma_to_ddr3_top_s1_waitrequest_from_sa;
  output           pb_dma_to_ddr3_top_s1_write;
  output  [ 31: 0] pb_dma_to_ddr3_top_s1_writedata;
  output           sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1;
  output           sgdma_rx_m_write_qualified_request_pb_dma_to_ddr3_top_s1;
  output           sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1;
  output           sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1;
  output           sgdma_tx_m_read_qualified_request_pb_dma_to_ddr3_top_s1;
  output           sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1;
  output           sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1_shift_register;
  output           sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1;
  input            clk;
  input            pb_dma_to_ddr3_top_s1_endofpacket;
  input   [ 31: 0] pb_dma_to_ddr3_top_s1_readdata;
  input            pb_dma_to_ddr3_top_s1_readdatavalid;
  input            pb_dma_to_ddr3_top_s1_waitrequest;
  input            reset_n;
  input   [ 31: 0] sgdma_rx_m_write_address_to_slave;
  input   [  3: 0] sgdma_rx_m_write_byteenable;
  input            sgdma_rx_m_write_write;
  input   [ 31: 0] sgdma_rx_m_write_writedata;
  input   [ 31: 0] sgdma_tx_m_read_address_to_slave;
  input            sgdma_tx_m_read_latency_counter;
  input            sgdma_tx_m_read_read;

  reg              d1_pb_dma_to_ddr3_top_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_pb_dma_to_ddr3_top_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_sgdma_rx_m_write_granted_slave_pb_dma_to_ddr3_top_s1;
  reg              last_cycle_sgdma_tx_m_read_granted_slave_pb_dma_to_ddr3_top_s1;
  wire    [ 24: 0] pb_dma_to_ddr3_top_s1_address;
  wire             pb_dma_to_ddr3_top_s1_allgrants;
  wire             pb_dma_to_ddr3_top_s1_allow_new_arb_cycle;
  wire             pb_dma_to_ddr3_top_s1_any_bursting_master_saved_grant;
  wire             pb_dma_to_ddr3_top_s1_any_continuerequest;
  reg     [  1: 0] pb_dma_to_ddr3_top_s1_arb_addend;
  wire             pb_dma_to_ddr3_top_s1_arb_counter_enable;
  reg     [  3: 0] pb_dma_to_ddr3_top_s1_arb_share_counter;
  wire    [  3: 0] pb_dma_to_ddr3_top_s1_arb_share_counter_next_value;
  wire    [  3: 0] pb_dma_to_ddr3_top_s1_arb_share_set_values;
  wire    [  1: 0] pb_dma_to_ddr3_top_s1_arb_winner;
  wire             pb_dma_to_ddr3_top_s1_arbiterlock;
  wire             pb_dma_to_ddr3_top_s1_arbiterlock2;
  wire             pb_dma_to_ddr3_top_s1_arbitration_holdoff_internal;
  wire             pb_dma_to_ddr3_top_s1_beginbursttransfer_internal;
  wire             pb_dma_to_ddr3_top_s1_begins_xfer;
  wire             pb_dma_to_ddr3_top_s1_burstcount;
  wire    [  3: 0] pb_dma_to_ddr3_top_s1_byteenable;
  wire             pb_dma_to_ddr3_top_s1_chipselect;
  wire    [  3: 0] pb_dma_to_ddr3_top_s1_chosen_master_double_vector;
  wire    [  1: 0] pb_dma_to_ddr3_top_s1_chosen_master_rot_left;
  wire             pb_dma_to_ddr3_top_s1_debugaccess;
  wire             pb_dma_to_ddr3_top_s1_end_xfer;
  wire             pb_dma_to_ddr3_top_s1_endofpacket_from_sa;
  wire             pb_dma_to_ddr3_top_s1_firsttransfer;
  wire    [  1: 0] pb_dma_to_ddr3_top_s1_grant_vector;
  wire             pb_dma_to_ddr3_top_s1_in_a_read_cycle;
  wire             pb_dma_to_ddr3_top_s1_in_a_write_cycle;
  wire    [  1: 0] pb_dma_to_ddr3_top_s1_master_qreq_vector;
  wire             pb_dma_to_ddr3_top_s1_move_on_to_next_transaction;
  wire    [ 24: 0] pb_dma_to_ddr3_top_s1_nativeaddress;
  wire             pb_dma_to_ddr3_top_s1_non_bursting_master_requests;
  wire             pb_dma_to_ddr3_top_s1_read;
  wire    [ 31: 0] pb_dma_to_ddr3_top_s1_readdata_from_sa;
  wire             pb_dma_to_ddr3_top_s1_readdatavalid_from_sa;
  reg              pb_dma_to_ddr3_top_s1_reg_firsttransfer;
  wire             pb_dma_to_ddr3_top_s1_reset_n;
  reg     [  1: 0] pb_dma_to_ddr3_top_s1_saved_chosen_master_vector;
  reg              pb_dma_to_ddr3_top_s1_slavearbiterlockenable;
  wire             pb_dma_to_ddr3_top_s1_slavearbiterlockenable2;
  wire             pb_dma_to_ddr3_top_s1_unreg_firsttransfer;
  wire             pb_dma_to_ddr3_top_s1_waitrequest_from_sa;
  wire             pb_dma_to_ddr3_top_s1_waits_for_read;
  wire             pb_dma_to_ddr3_top_s1_waits_for_write;
  wire             pb_dma_to_ddr3_top_s1_write;
  wire    [ 31: 0] pb_dma_to_ddr3_top_s1_writedata;
  wire             sgdma_rx_m_write_arbiterlock;
  wire             sgdma_rx_m_write_arbiterlock2;
  wire             sgdma_rx_m_write_continuerequest;
  wire             sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1;
  wire             sgdma_rx_m_write_qualified_request_pb_dma_to_ddr3_top_s1;
  wire             sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1;
  wire             sgdma_rx_m_write_saved_grant_pb_dma_to_ddr3_top_s1;
  wire             sgdma_tx_m_read_arbiterlock;
  wire             sgdma_tx_m_read_arbiterlock2;
  wire             sgdma_tx_m_read_continuerequest;
  wire             sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1;
  wire             sgdma_tx_m_read_qualified_request_pb_dma_to_ddr3_top_s1;
  wire             sgdma_tx_m_read_rdv_fifo_empty_pb_dma_to_ddr3_top_s1;
  wire             sgdma_tx_m_read_rdv_fifo_output_from_pb_dma_to_ddr3_top_s1;
  wire             sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1;
  wire             sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1_shift_register;
  wire             sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1;
  wire             sgdma_tx_m_read_saved_grant_pb_dma_to_ddr3_top_s1;
  wire    [ 31: 0] shifted_address_to_pb_dma_to_ddr3_top_s1_from_sgdma_rx_m_write;
  wire    [ 31: 0] shifted_address_to_pb_dma_to_ddr3_top_s1_from_sgdma_tx_m_read;
  wire             wait_for_pb_dma_to_ddr3_top_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~pb_dma_to_ddr3_top_s1_end_xfer;
    end


  assign pb_dma_to_ddr3_top_s1_begins_xfer = ~d1_reasons_to_wait & ((sgdma_rx_m_write_qualified_request_pb_dma_to_ddr3_top_s1 | sgdma_tx_m_read_qualified_request_pb_dma_to_ddr3_top_s1));
  //assign pb_dma_to_ddr3_top_s1_readdata_from_sa = pb_dma_to_ddr3_top_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_readdata_from_sa = pb_dma_to_ddr3_top_s1_readdata;

  assign sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1 = (({sgdma_rx_m_write_address_to_slave[31 : 27] , 27'b0} == 32'h10000000) & (sgdma_rx_m_write_write)) & sgdma_rx_m_write_write;
  //assign pb_dma_to_ddr3_top_s1_waitrequest_from_sa = pb_dma_to_ddr3_top_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_waitrequest_from_sa = pb_dma_to_ddr3_top_s1_waitrequest;

  //pb_dma_to_ddr3_top_s1_arb_share_counter set values, which is an e_mux
  assign pb_dma_to_ddr3_top_s1_arb_share_set_values = (sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1)? 8 :
    (sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1)? 8 :
    (sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1)? 8 :
    (sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1)? 8 :
    (sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1)? 8 :
    (sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1)? 8 :
    1;

  //pb_dma_to_ddr3_top_s1_non_bursting_master_requests mux, which is an e_mux
  assign pb_dma_to_ddr3_top_s1_non_bursting_master_requests = sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1 |
    sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1 |
    sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1 |
    sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1 |
    sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1 |
    sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1;

  //pb_dma_to_ddr3_top_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign pb_dma_to_ddr3_top_s1_any_bursting_master_saved_grant = 0;

  //pb_dma_to_ddr3_top_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_arb_share_counter_next_value = pb_dma_to_ddr3_top_s1_firsttransfer ? (pb_dma_to_ddr3_top_s1_arb_share_set_values - 1) : |pb_dma_to_ddr3_top_s1_arb_share_counter ? (pb_dma_to_ddr3_top_s1_arb_share_counter - 1) : 0;

  //pb_dma_to_ddr3_top_s1_allgrants all slave grants, which is an e_mux
  assign pb_dma_to_ddr3_top_s1_allgrants = (|pb_dma_to_ddr3_top_s1_grant_vector) |
    (|pb_dma_to_ddr3_top_s1_grant_vector) |
    (|pb_dma_to_ddr3_top_s1_grant_vector) |
    (|pb_dma_to_ddr3_top_s1_grant_vector) |
    (|pb_dma_to_ddr3_top_s1_grant_vector) |
    (|pb_dma_to_ddr3_top_s1_grant_vector);

  //pb_dma_to_ddr3_top_s1_end_xfer assignment, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_end_xfer = ~(pb_dma_to_ddr3_top_s1_waits_for_read | pb_dma_to_ddr3_top_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_pb_dma_to_ddr3_top_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_pb_dma_to_ddr3_top_s1 = pb_dma_to_ddr3_top_s1_end_xfer & (~pb_dma_to_ddr3_top_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //pb_dma_to_ddr3_top_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_pb_dma_to_ddr3_top_s1 & pb_dma_to_ddr3_top_s1_allgrants) | (end_xfer_arb_share_counter_term_pb_dma_to_ddr3_top_s1 & ~pb_dma_to_ddr3_top_s1_non_bursting_master_requests);

  //pb_dma_to_ddr3_top_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_ddr3_top_s1_arb_share_counter <= 0;
      else if (pb_dma_to_ddr3_top_s1_arb_counter_enable)
          pb_dma_to_ddr3_top_s1_arb_share_counter <= pb_dma_to_ddr3_top_s1_arb_share_counter_next_value;
    end


  //pb_dma_to_ddr3_top_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_ddr3_top_s1_slavearbiterlockenable <= 0;
      else if ((|pb_dma_to_ddr3_top_s1_master_qreq_vector & end_xfer_arb_share_counter_term_pb_dma_to_ddr3_top_s1) | (end_xfer_arb_share_counter_term_pb_dma_to_ddr3_top_s1 & ~pb_dma_to_ddr3_top_s1_non_bursting_master_requests))
          pb_dma_to_ddr3_top_s1_slavearbiterlockenable <= |pb_dma_to_ddr3_top_s1_arb_share_counter_next_value;
    end


  //sgdma_rx/m_write pb_dma_to_ddr3_top/s1 arbiterlock, which is an e_assign
  assign sgdma_rx_m_write_arbiterlock = pb_dma_to_ddr3_top_s1_slavearbiterlockenable & sgdma_rx_m_write_continuerequest;

  //pb_dma_to_ddr3_top_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_slavearbiterlockenable2 = |pb_dma_to_ddr3_top_s1_arb_share_counter_next_value;

  //sgdma_rx/m_write pb_dma_to_ddr3_top/s1 arbiterlock2, which is an e_assign
  assign sgdma_rx_m_write_arbiterlock2 = pb_dma_to_ddr3_top_s1_slavearbiterlockenable2 & sgdma_rx_m_write_continuerequest;

  //sgdma_tx/m_read pb_dma_to_ddr3_top/s1 arbiterlock, which is an e_assign
  assign sgdma_tx_m_read_arbiterlock = pb_dma_to_ddr3_top_s1_slavearbiterlockenable & sgdma_tx_m_read_continuerequest;

  //sgdma_tx/m_read pb_dma_to_ddr3_top/s1 arbiterlock2, which is an e_assign
  assign sgdma_tx_m_read_arbiterlock2 = pb_dma_to_ddr3_top_s1_slavearbiterlockenable2 & sgdma_tx_m_read_continuerequest;

  //sgdma_tx/m_read granted pb_dma_to_ddr3_top/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_tx_m_read_granted_slave_pb_dma_to_ddr3_top_s1 <= 0;
      else 
        last_cycle_sgdma_tx_m_read_granted_slave_pb_dma_to_ddr3_top_s1 <= sgdma_tx_m_read_saved_grant_pb_dma_to_ddr3_top_s1 ? 1 : (pb_dma_to_ddr3_top_s1_arbitration_holdoff_internal | ~sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1) ? 0 : last_cycle_sgdma_tx_m_read_granted_slave_pb_dma_to_ddr3_top_s1;
    end


  //sgdma_tx_m_read_continuerequest continued request, which is an e_mux
  assign sgdma_tx_m_read_continuerequest = last_cycle_sgdma_tx_m_read_granted_slave_pb_dma_to_ddr3_top_s1 & sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1;

  //pb_dma_to_ddr3_top_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign pb_dma_to_ddr3_top_s1_any_continuerequest = sgdma_tx_m_read_continuerequest |
    sgdma_rx_m_write_continuerequest;

  assign sgdma_rx_m_write_qualified_request_pb_dma_to_ddr3_top_s1 = sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1 & ~(sgdma_tx_m_read_arbiterlock);
  //pb_dma_to_ddr3_top_s1_writedata mux, which is an e_mux
  assign pb_dma_to_ddr3_top_s1_writedata = sgdma_rx_m_write_writedata;

  //assign pb_dma_to_ddr3_top_s1_endofpacket_from_sa = pb_dma_to_ddr3_top_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_endofpacket_from_sa = pb_dma_to_ddr3_top_s1_endofpacket;

  assign sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1 = (({sgdma_tx_m_read_address_to_slave[31 : 27] , 27'b0} == 32'h10000000) & (sgdma_tx_m_read_read)) & sgdma_tx_m_read_read;
  //assign pb_dma_to_ddr3_top_s1_readdatavalid_from_sa = pb_dma_to_ddr3_top_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_readdatavalid_from_sa = pb_dma_to_ddr3_top_s1_readdatavalid;

  //sgdma_rx/m_write granted pb_dma_to_ddr3_top/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_rx_m_write_granted_slave_pb_dma_to_ddr3_top_s1 <= 0;
      else 
        last_cycle_sgdma_rx_m_write_granted_slave_pb_dma_to_ddr3_top_s1 <= sgdma_rx_m_write_saved_grant_pb_dma_to_ddr3_top_s1 ? 1 : (pb_dma_to_ddr3_top_s1_arbitration_holdoff_internal | ~sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1) ? 0 : last_cycle_sgdma_rx_m_write_granted_slave_pb_dma_to_ddr3_top_s1;
    end


  //sgdma_rx_m_write_continuerequest continued request, which is an e_mux
  assign sgdma_rx_m_write_continuerequest = last_cycle_sgdma_rx_m_write_granted_slave_pb_dma_to_ddr3_top_s1 & sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1;

  assign sgdma_tx_m_read_qualified_request_pb_dma_to_ddr3_top_s1 = sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1 & ~((sgdma_tx_m_read_read & ((sgdma_tx_m_read_latency_counter != 0) | (1 < sgdma_tx_m_read_latency_counter))) | sgdma_rx_m_write_arbiterlock);
  //unique name for pb_dma_to_ddr3_top_s1_move_on_to_next_transaction, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_move_on_to_next_transaction = pb_dma_to_ddr3_top_s1_readdatavalid_from_sa;

  //rdv_fifo_for_sgdma_tx_m_read_to_pb_dma_to_ddr3_top_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_sgdma_tx_m_read_to_pb_dma_to_ddr3_top_s1_module rdv_fifo_for_sgdma_tx_m_read_to_pb_dma_to_ddr3_top_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1),
      .data_out             (sgdma_tx_m_read_rdv_fifo_output_from_pb_dma_to_ddr3_top_s1),
      .empty                (),
      .fifo_contains_ones_n (sgdma_tx_m_read_rdv_fifo_empty_pb_dma_to_ddr3_top_s1),
      .full                 (),
      .read                 (pb_dma_to_ddr3_top_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~pb_dma_to_ddr3_top_s1_waits_for_read)
    );

  assign sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1_shift_register = ~sgdma_tx_m_read_rdv_fifo_empty_pb_dma_to_ddr3_top_s1;
  //local readdatavalid sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1, which is an e_mux
  assign sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1 = (pb_dma_to_ddr3_top_s1_readdatavalid_from_sa & sgdma_tx_m_read_rdv_fifo_output_from_pb_dma_to_ddr3_top_s1) & ~ sgdma_tx_m_read_rdv_fifo_empty_pb_dma_to_ddr3_top_s1;

  //allow new arb cycle for pb_dma_to_ddr3_top/s1, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_allow_new_arb_cycle = ~sgdma_rx_m_write_arbiterlock & ~sgdma_tx_m_read_arbiterlock;

  //sgdma_tx/m_read assignment into master qualified-requests vector for pb_dma_to_ddr3_top/s1, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_master_qreq_vector[0] = sgdma_tx_m_read_qualified_request_pb_dma_to_ddr3_top_s1;

  //sgdma_tx/m_read grant pb_dma_to_ddr3_top/s1, which is an e_assign
  assign sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1 = pb_dma_to_ddr3_top_s1_grant_vector[0];

  //sgdma_tx/m_read saved-grant pb_dma_to_ddr3_top/s1, which is an e_assign
  assign sgdma_tx_m_read_saved_grant_pb_dma_to_ddr3_top_s1 = pb_dma_to_ddr3_top_s1_arb_winner[0] && sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1;

  //sgdma_rx/m_write assignment into master qualified-requests vector for pb_dma_to_ddr3_top/s1, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_master_qreq_vector[1] = sgdma_rx_m_write_qualified_request_pb_dma_to_ddr3_top_s1;

  //sgdma_rx/m_write grant pb_dma_to_ddr3_top/s1, which is an e_assign
  assign sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1 = pb_dma_to_ddr3_top_s1_grant_vector[1];

  //sgdma_rx/m_write saved-grant pb_dma_to_ddr3_top/s1, which is an e_assign
  assign sgdma_rx_m_write_saved_grant_pb_dma_to_ddr3_top_s1 = pb_dma_to_ddr3_top_s1_arb_winner[1] && sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1;

  //pb_dma_to_ddr3_top/s1 chosen-master double-vector, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_chosen_master_double_vector = {pb_dma_to_ddr3_top_s1_master_qreq_vector, pb_dma_to_ddr3_top_s1_master_qreq_vector} & ({~pb_dma_to_ddr3_top_s1_master_qreq_vector, ~pb_dma_to_ddr3_top_s1_master_qreq_vector} + pb_dma_to_ddr3_top_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign pb_dma_to_ddr3_top_s1_arb_winner = (pb_dma_to_ddr3_top_s1_allow_new_arb_cycle & | pb_dma_to_ddr3_top_s1_grant_vector) ? pb_dma_to_ddr3_top_s1_grant_vector : pb_dma_to_ddr3_top_s1_saved_chosen_master_vector;

  //saved pb_dma_to_ddr3_top_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_ddr3_top_s1_saved_chosen_master_vector <= 0;
      else if (pb_dma_to_ddr3_top_s1_allow_new_arb_cycle)
          pb_dma_to_ddr3_top_s1_saved_chosen_master_vector <= |pb_dma_to_ddr3_top_s1_grant_vector ? pb_dma_to_ddr3_top_s1_grant_vector : pb_dma_to_ddr3_top_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign pb_dma_to_ddr3_top_s1_grant_vector = {(pb_dma_to_ddr3_top_s1_chosen_master_double_vector[1] | pb_dma_to_ddr3_top_s1_chosen_master_double_vector[3]),
    (pb_dma_to_ddr3_top_s1_chosen_master_double_vector[0] | pb_dma_to_ddr3_top_s1_chosen_master_double_vector[2])};

  //pb_dma_to_ddr3_top/s1 chosen master rotated left, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_chosen_master_rot_left = (pb_dma_to_ddr3_top_s1_arb_winner << 1) ? (pb_dma_to_ddr3_top_s1_arb_winner << 1) : 1;

  //pb_dma_to_ddr3_top/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_ddr3_top_s1_arb_addend <= 1;
      else if (|pb_dma_to_ddr3_top_s1_grant_vector)
          pb_dma_to_ddr3_top_s1_arb_addend <= pb_dma_to_ddr3_top_s1_end_xfer? pb_dma_to_ddr3_top_s1_chosen_master_rot_left : pb_dma_to_ddr3_top_s1_grant_vector;
    end


  //pb_dma_to_ddr3_top_s1_reset_n assignment, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_reset_n = reset_n;

  assign pb_dma_to_ddr3_top_s1_chipselect = sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1 | sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1;
  //pb_dma_to_ddr3_top_s1_firsttransfer first transaction, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_firsttransfer = pb_dma_to_ddr3_top_s1_begins_xfer ? pb_dma_to_ddr3_top_s1_unreg_firsttransfer : pb_dma_to_ddr3_top_s1_reg_firsttransfer;

  //pb_dma_to_ddr3_top_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_unreg_firsttransfer = ~(pb_dma_to_ddr3_top_s1_slavearbiterlockenable & pb_dma_to_ddr3_top_s1_any_continuerequest);

  //pb_dma_to_ddr3_top_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_ddr3_top_s1_reg_firsttransfer <= 1'b1;
      else if (pb_dma_to_ddr3_top_s1_begins_xfer)
          pb_dma_to_ddr3_top_s1_reg_firsttransfer <= pb_dma_to_ddr3_top_s1_unreg_firsttransfer;
    end


  //pb_dma_to_ddr3_top_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_beginbursttransfer_internal = pb_dma_to_ddr3_top_s1_begins_xfer;

  //pb_dma_to_ddr3_top_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_arbitration_holdoff_internal = pb_dma_to_ddr3_top_s1_begins_xfer & pb_dma_to_ddr3_top_s1_firsttransfer;

  //pb_dma_to_ddr3_top_s1_read assignment, which is an e_mux
  assign pb_dma_to_ddr3_top_s1_read = sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1 & sgdma_tx_m_read_read;

  //pb_dma_to_ddr3_top_s1_write assignment, which is an e_mux
  assign pb_dma_to_ddr3_top_s1_write = sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1 & sgdma_rx_m_write_write;

  assign shifted_address_to_pb_dma_to_ddr3_top_s1_from_sgdma_rx_m_write = sgdma_rx_m_write_address_to_slave;
  //pb_dma_to_ddr3_top_s1_address mux, which is an e_mux
  assign pb_dma_to_ddr3_top_s1_address = (sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1)? (shifted_address_to_pb_dma_to_ddr3_top_s1_from_sgdma_rx_m_write >> 2) :
    (shifted_address_to_pb_dma_to_ddr3_top_s1_from_sgdma_tx_m_read >> 2);

  assign shifted_address_to_pb_dma_to_ddr3_top_s1_from_sgdma_tx_m_read = sgdma_tx_m_read_address_to_slave;
  //slaveid pb_dma_to_ddr3_top_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign pb_dma_to_ddr3_top_s1_nativeaddress = (sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1)? (sgdma_rx_m_write_address_to_slave >> 2) :
    (sgdma_tx_m_read_address_to_slave >> 2);

  //d1_pb_dma_to_ddr3_top_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_pb_dma_to_ddr3_top_s1_end_xfer <= 1;
      else 
        d1_pb_dma_to_ddr3_top_s1_end_xfer <= pb_dma_to_ddr3_top_s1_end_xfer;
    end


  //pb_dma_to_ddr3_top_s1_waits_for_read in a cycle, which is an e_mux
  assign pb_dma_to_ddr3_top_s1_waits_for_read = pb_dma_to_ddr3_top_s1_in_a_read_cycle & pb_dma_to_ddr3_top_s1_waitrequest_from_sa;

  //pb_dma_to_ddr3_top_s1_in_a_read_cycle assignment, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_in_a_read_cycle = sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1 & sgdma_tx_m_read_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = pb_dma_to_ddr3_top_s1_in_a_read_cycle;

  //pb_dma_to_ddr3_top_s1_waits_for_write in a cycle, which is an e_mux
  assign pb_dma_to_ddr3_top_s1_waits_for_write = pb_dma_to_ddr3_top_s1_in_a_write_cycle & pb_dma_to_ddr3_top_s1_waitrequest_from_sa;

  //pb_dma_to_ddr3_top_s1_in_a_write_cycle assignment, which is an e_assign
  assign pb_dma_to_ddr3_top_s1_in_a_write_cycle = sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1 & sgdma_rx_m_write_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = pb_dma_to_ddr3_top_s1_in_a_write_cycle;

  assign wait_for_pb_dma_to_ddr3_top_s1_counter = 0;
  //pb_dma_to_ddr3_top_s1_byteenable byte enable port mux, which is an e_mux
  assign pb_dma_to_ddr3_top_s1_byteenable = (sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1)? sgdma_rx_m_write_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign pb_dma_to_ddr3_top_s1_burstcount = 1;

  //pb_dma_to_ddr3_top/s1 arbiterlock assigned from _handle_arbiterlock, which is an e_mux
  assign pb_dma_to_ddr3_top_s1_arbiterlock = (sgdma_rx_m_write_arbiterlock)? sgdma_rx_m_write_arbiterlock :
    sgdma_tx_m_read_arbiterlock;

  //pb_dma_to_ddr3_top/s1 arbiterlock2 assigned from _handle_arbiterlock2, which is an e_mux
  assign pb_dma_to_ddr3_top_s1_arbiterlock2 = (sgdma_rx_m_write_arbiterlock2)? sgdma_rx_m_write_arbiterlock2 :
    sgdma_tx_m_read_arbiterlock2;

  //debugaccess mux, which is an e_mux
  assign pb_dma_to_ddr3_top_s1_debugaccess = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pb_dma_to_ddr3_top/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1 + sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (sgdma_rx_m_write_saved_grant_pb_dma_to_ddr3_top_s1 + sgdma_tx_m_read_saved_grant_pb_dma_to_ddr3_top_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo_module (
                                                                      // inputs:
                                                                       clear_fifo,
                                                                       clk,
                                                                       data_in,
                                                                       read,
                                                                       reset_n,
                                                                       sync_reset,
                                                                       write,

                                                                      // outputs:
                                                                       data_out,
                                                                       empty,
                                                                       fifo_contains_ones_n,
                                                                       full
                                                                    )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  wire             full_32;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_31;
  assign empty = !full_0;
  assign full_32 = 0;
  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    0;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pb_dma_to_ddr3_top_m1_arbitrator (
                                          // inputs:
                                           clk,
                                           d1_ddr3_top_s1_end_xfer,
                                           ddr3_top_s1_readdata_from_sa,
                                           ddr3_top_s1_waitrequest_n_from_sa,
                                           pb_dma_to_ddr3_top_m1_address,
                                           pb_dma_to_ddr3_top_m1_burstcount,
                                           pb_dma_to_ddr3_top_m1_byteenable,
                                           pb_dma_to_ddr3_top_m1_chipselect,
                                           pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1,
                                           pb_dma_to_ddr3_top_m1_qualified_request_ddr3_top_s1,
                                           pb_dma_to_ddr3_top_m1_read,
                                           pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1,
                                           pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register,
                                           pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1,
                                           pb_dma_to_ddr3_top_m1_write,
                                           pb_dma_to_ddr3_top_m1_writedata,
                                           reset_n,

                                          // outputs:
                                           pb_dma_to_ddr3_top_m1_address_to_slave,
                                           pb_dma_to_ddr3_top_m1_latency_counter,
                                           pb_dma_to_ddr3_top_m1_readdata,
                                           pb_dma_to_ddr3_top_m1_readdatavalid,
                                           pb_dma_to_ddr3_top_m1_waitrequest
                                        )
;

  output  [ 26: 0] pb_dma_to_ddr3_top_m1_address_to_slave;
  output           pb_dma_to_ddr3_top_m1_latency_counter;
  output  [ 31: 0] pb_dma_to_ddr3_top_m1_readdata;
  output           pb_dma_to_ddr3_top_m1_readdatavalid;
  output           pb_dma_to_ddr3_top_m1_waitrequest;
  input            clk;
  input            d1_ddr3_top_s1_end_xfer;
  input   [ 63: 0] ddr3_top_s1_readdata_from_sa;
  input            ddr3_top_s1_waitrequest_n_from_sa;
  input   [ 26: 0] pb_dma_to_ddr3_top_m1_address;
  input            pb_dma_to_ddr3_top_m1_burstcount;
  input   [  3: 0] pb_dma_to_ddr3_top_m1_byteenable;
  input            pb_dma_to_ddr3_top_m1_chipselect;
  input            pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1;
  input            pb_dma_to_ddr3_top_m1_qualified_request_ddr3_top_s1;
  input            pb_dma_to_ddr3_top_m1_read;
  input            pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1;
  input            pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register;
  input            pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1;
  input            pb_dma_to_ddr3_top_m1_write;
  input   [ 31: 0] pb_dma_to_ddr3_top_m1_writedata;
  input            reset_n;

  reg              active_and_waiting_last_time;
  wire    [ 31: 0] ddr3_top_s1_readdata_from_sa_part_selected_by_negative_dbs;
  wire             empty_selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo;
  wire             full_selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo;
  wire             latency_load_value;
  wire             p1_pb_dma_to_ddr3_top_m1_latency_counter;
  reg     [ 26: 0] pb_dma_to_ddr3_top_m1_address_last_time;
  wire    [ 26: 0] pb_dma_to_ddr3_top_m1_address_to_slave;
  reg              pb_dma_to_ddr3_top_m1_burstcount_last_time;
  reg     [  3: 0] pb_dma_to_ddr3_top_m1_byteenable_last_time;
  reg              pb_dma_to_ddr3_top_m1_chipselect_last_time;
  wire             pb_dma_to_ddr3_top_m1_is_granted_some_slave;
  reg              pb_dma_to_ddr3_top_m1_latency_counter;
  reg              pb_dma_to_ddr3_top_m1_read_but_no_slave_selected;
  reg              pb_dma_to_ddr3_top_m1_read_last_time;
  wire    [ 31: 0] pb_dma_to_ddr3_top_m1_readdata;
  wire             pb_dma_to_ddr3_top_m1_readdatavalid;
  wire             pb_dma_to_ddr3_top_m1_run;
  wire             pb_dma_to_ddr3_top_m1_waitrequest;
  reg              pb_dma_to_ddr3_top_m1_write_last_time;
  reg     [ 31: 0] pb_dma_to_ddr3_top_m1_writedata_last_time;
  wire             pre_flush_pb_dma_to_ddr3_top_m1_readdatavalid;
  wire             r_0;
  wire             read_selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo;
  wire             selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo_output;
  wire             selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo_output_ddr3_top_s1;
  wire             write_selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (pb_dma_to_ddr3_top_m1_qualified_request_ddr3_top_s1 | ~pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1) & (pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1 | ~pb_dma_to_ddr3_top_m1_qualified_request_ddr3_top_s1) & ((~pb_dma_to_ddr3_top_m1_qualified_request_ddr3_top_s1 | ~pb_dma_to_ddr3_top_m1_chipselect | (1 & ddr3_top_s1_waitrequest_n_from_sa & pb_dma_to_ddr3_top_m1_chipselect))) & ((~pb_dma_to_ddr3_top_m1_qualified_request_ddr3_top_s1 | ~pb_dma_to_ddr3_top_m1_chipselect | (1 & ddr3_top_s1_waitrequest_n_from_sa & pb_dma_to_ddr3_top_m1_chipselect)));

  //cascaded wait assignment, which is an e_assign
  assign pb_dma_to_ddr3_top_m1_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign pb_dma_to_ddr3_top_m1_address_to_slave = pb_dma_to_ddr3_top_m1_address[26 : 0];

  //pb_dma_to_ddr3_top_m1_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_ddr3_top_m1_read_but_no_slave_selected <= 0;
      else 
        pb_dma_to_ddr3_top_m1_read_but_no_slave_selected <= (pb_dma_to_ddr3_top_m1_read & pb_dma_to_ddr3_top_m1_chipselect) & pb_dma_to_ddr3_top_m1_run & ~pb_dma_to_ddr3_top_m1_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign pb_dma_to_ddr3_top_m1_is_granted_some_slave = pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_pb_dma_to_ddr3_top_m1_readdatavalid = pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign pb_dma_to_ddr3_top_m1_readdatavalid = pb_dma_to_ddr3_top_m1_read_but_no_slave_selected |
    pre_flush_pb_dma_to_ddr3_top_m1_readdatavalid;

  //Negative Dynamic Bus-sizing mux.
  //this mux selects the correct half of the 
  //wide data coming from the slave ddr3_top/s1 
  assign ddr3_top_s1_readdata_from_sa_part_selected_by_negative_dbs = ((selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo_output_ddr3_top_s1 == 0))? ddr3_top_s1_readdata_from_sa[31 : 0] :
    ddr3_top_s1_readdata_from_sa[63 : 32];

  //read_selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo fifo read, which is an e_mux
  assign read_selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo = pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1;

  //write_selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo fifo write, which is an e_mux
  assign write_selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo = (pb_dma_to_ddr3_top_m1_read & pb_dma_to_ddr3_top_m1_chipselect) & pb_dma_to_ddr3_top_m1_run & pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1;

  assign selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo_output_ddr3_top_s1 = selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo_output;
  //selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo, which is an e_fifo_with_registered_outputs
  selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo_module selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (pb_dma_to_ddr3_top_m1_address_to_slave[2]),
      .data_out             (selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo_output),
      .empty                (empty_selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo),
      .fifo_contains_ones_n (),
      .full                 (full_selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo),
      .read                 (read_selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (write_selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo)
    );

  //pb_dma_to_ddr3_top/m1 readdata mux, which is an e_mux
  assign pb_dma_to_ddr3_top_m1_readdata = ddr3_top_s1_readdata_from_sa_part_selected_by_negative_dbs;

  //actual waitrequest port, which is an e_assign
  assign pb_dma_to_ddr3_top_m1_waitrequest = ~pb_dma_to_ddr3_top_m1_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_ddr3_top_m1_latency_counter <= 0;
      else 
        pb_dma_to_ddr3_top_m1_latency_counter <= p1_pb_dma_to_ddr3_top_m1_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_pb_dma_to_ddr3_top_m1_latency_counter = ((pb_dma_to_ddr3_top_m1_run & (pb_dma_to_ddr3_top_m1_read & pb_dma_to_ddr3_top_m1_chipselect)))? latency_load_value :
    (pb_dma_to_ddr3_top_m1_latency_counter)? pb_dma_to_ddr3_top_m1_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pb_dma_to_ddr3_top_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_ddr3_top_m1_address_last_time <= 0;
      else 
        pb_dma_to_ddr3_top_m1_address_last_time <= pb_dma_to_ddr3_top_m1_address;
    end


  //pb_dma_to_ddr3_top/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= pb_dma_to_ddr3_top_m1_waitrequest & pb_dma_to_ddr3_top_m1_chipselect;
    end


  //pb_dma_to_ddr3_top_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_dma_to_ddr3_top_m1_address != pb_dma_to_ddr3_top_m1_address_last_time))
        begin
          $write("%0d ns: pb_dma_to_ddr3_top_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_dma_to_ddr3_top_m1_chipselect check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_ddr3_top_m1_chipselect_last_time <= 0;
      else 
        pb_dma_to_ddr3_top_m1_chipselect_last_time <= pb_dma_to_ddr3_top_m1_chipselect;
    end


  //pb_dma_to_ddr3_top_m1_chipselect matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_dma_to_ddr3_top_m1_chipselect != pb_dma_to_ddr3_top_m1_chipselect_last_time))
        begin
          $write("%0d ns: pb_dma_to_ddr3_top_m1_chipselect did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_dma_to_ddr3_top_m1_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_ddr3_top_m1_burstcount_last_time <= 0;
      else 
        pb_dma_to_ddr3_top_m1_burstcount_last_time <= pb_dma_to_ddr3_top_m1_burstcount;
    end


  //pb_dma_to_ddr3_top_m1_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_dma_to_ddr3_top_m1_burstcount != pb_dma_to_ddr3_top_m1_burstcount_last_time))
        begin
          $write("%0d ns: pb_dma_to_ddr3_top_m1_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_dma_to_ddr3_top_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_ddr3_top_m1_byteenable_last_time <= 0;
      else 
        pb_dma_to_ddr3_top_m1_byteenable_last_time <= pb_dma_to_ddr3_top_m1_byteenable;
    end


  //pb_dma_to_ddr3_top_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_dma_to_ddr3_top_m1_byteenable != pb_dma_to_ddr3_top_m1_byteenable_last_time))
        begin
          $write("%0d ns: pb_dma_to_ddr3_top_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_dma_to_ddr3_top_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_ddr3_top_m1_read_last_time <= 0;
      else 
        pb_dma_to_ddr3_top_m1_read_last_time <= pb_dma_to_ddr3_top_m1_read;
    end


  //pb_dma_to_ddr3_top_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_dma_to_ddr3_top_m1_read != pb_dma_to_ddr3_top_m1_read_last_time))
        begin
          $write("%0d ns: pb_dma_to_ddr3_top_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_dma_to_ddr3_top_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_ddr3_top_m1_write_last_time <= 0;
      else 
        pb_dma_to_ddr3_top_m1_write_last_time <= pb_dma_to_ddr3_top_m1_write;
    end


  //pb_dma_to_ddr3_top_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_dma_to_ddr3_top_m1_write != pb_dma_to_ddr3_top_m1_write_last_time))
        begin
          $write("%0d ns: pb_dma_to_ddr3_top_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_dma_to_ddr3_top_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_ddr3_top_m1_writedata_last_time <= 0;
      else 
        pb_dma_to_ddr3_top_m1_writedata_last_time <= pb_dma_to_ddr3_top_m1_writedata;
    end


  //pb_dma_to_ddr3_top_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_dma_to_ddr3_top_m1_writedata != pb_dma_to_ddr3_top_m1_writedata_last_time) & (pb_dma_to_ddr3_top_m1_write & pb_dma_to_ddr3_top_m1_chipselect))
        begin
          $write("%0d ns: pb_dma_to_ddr3_top_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end


  //selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo read when empty, which is an e_process
  always @(posedge clk)
    begin
      if (empty_selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo & read_selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo)
        begin
          $write("%0d ns: pb_dma_to_ddr3_top/m1 negative rdv fifo selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo: read AND empty.\n", $time);
          $stop;
        end
    end


  //selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo write when full, which is an e_process
  always @(posedge clk)
    begin
      if (full_selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo & write_selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo & ~read_selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo)
        begin
          $write("%0d ns: pb_dma_to_ddr3_top/m1 negative rdv fifo selecto_nrdv_pb_dma_to_ddr3_top_m1_1_ddr3_top_s1_fifo: write AND full.\n", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pb_dma_to_ddr3_top_bridge_arbitrator 
;



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_sgdma_rx_descriptor_read_to_pb_dma_to_descriptor_memory_s1_module (
                                                                                        // inputs:
                                                                                         clear_fifo,
                                                                                         clk,
                                                                                         data_in,
                                                                                         read,
                                                                                         reset_n,
                                                                                         sync_reset,
                                                                                         write,

                                                                                        // outputs:
                                                                                         data_out,
                                                                                         empty,
                                                                                         fifo_contains_ones_n,
                                                                                         full
                                                                                      )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_sgdma_tx_descriptor_read_to_pb_dma_to_descriptor_memory_s1_module (
                                                                                        // inputs:
                                                                                         clear_fifo,
                                                                                         clk,
                                                                                         data_in,
                                                                                         read,
                                                                                         reset_n,
                                                                                         sync_reset,
                                                                                         write,

                                                                                        // outputs:
                                                                                         data_out,
                                                                                         empty,
                                                                                         fifo_contains_ones_n,
                                                                                         full
                                                                                      )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pb_dma_to_descriptor_memory_s1_arbitrator (
                                                   // inputs:
                                                    clk,
                                                    pb_dma_to_descriptor_memory_s1_endofpacket,
                                                    pb_dma_to_descriptor_memory_s1_readdata,
                                                    pb_dma_to_descriptor_memory_s1_readdatavalid,
                                                    pb_dma_to_descriptor_memory_s1_waitrequest,
                                                    reset_n,
                                                    sgdma_rx_descriptor_read_address_to_slave,
                                                    sgdma_rx_descriptor_read_latency_counter,
                                                    sgdma_rx_descriptor_read_read,
                                                    sgdma_rx_descriptor_write_address_to_slave,
                                                    sgdma_rx_descriptor_write_write,
                                                    sgdma_rx_descriptor_write_writedata,
                                                    sgdma_tx_descriptor_read_address_to_slave,
                                                    sgdma_tx_descriptor_read_latency_counter,
                                                    sgdma_tx_descriptor_read_read,
                                                    sgdma_tx_descriptor_write_address_to_slave,
                                                    sgdma_tx_descriptor_write_write,
                                                    sgdma_tx_descriptor_write_writedata,

                                                   // outputs:
                                                    d1_pb_dma_to_descriptor_memory_s1_end_xfer,
                                                    pb_dma_to_descriptor_memory_s1_address,
                                                    pb_dma_to_descriptor_memory_s1_arbiterlock,
                                                    pb_dma_to_descriptor_memory_s1_arbiterlock2,
                                                    pb_dma_to_descriptor_memory_s1_burstcount,
                                                    pb_dma_to_descriptor_memory_s1_byteenable,
                                                    pb_dma_to_descriptor_memory_s1_chipselect,
                                                    pb_dma_to_descriptor_memory_s1_debugaccess,
                                                    pb_dma_to_descriptor_memory_s1_endofpacket_from_sa,
                                                    pb_dma_to_descriptor_memory_s1_nativeaddress,
                                                    pb_dma_to_descriptor_memory_s1_read,
                                                    pb_dma_to_descriptor_memory_s1_readdata_from_sa,
                                                    pb_dma_to_descriptor_memory_s1_reset_n,
                                                    pb_dma_to_descriptor_memory_s1_waitrequest_from_sa,
                                                    pb_dma_to_descriptor_memory_s1_write,
                                                    pb_dma_to_descriptor_memory_s1_writedata,
                                                    sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1,
                                                    sgdma_rx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1,
                                                    sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1,
                                                    sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register,
                                                    sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1,
                                                    sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1,
                                                    sgdma_rx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1,
                                                    sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1,
                                                    sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1,
                                                    sgdma_tx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1,
                                                    sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1,
                                                    sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register,
                                                    sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1,
                                                    sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1,
                                                    sgdma_tx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1,
                                                    sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1
                                                 )
;

  output           d1_pb_dma_to_descriptor_memory_s1_end_xfer;
  output  [ 11: 0] pb_dma_to_descriptor_memory_s1_address;
  output           pb_dma_to_descriptor_memory_s1_arbiterlock;
  output           pb_dma_to_descriptor_memory_s1_arbiterlock2;
  output           pb_dma_to_descriptor_memory_s1_burstcount;
  output  [  3: 0] pb_dma_to_descriptor_memory_s1_byteenable;
  output           pb_dma_to_descriptor_memory_s1_chipselect;
  output           pb_dma_to_descriptor_memory_s1_debugaccess;
  output           pb_dma_to_descriptor_memory_s1_endofpacket_from_sa;
  output  [ 11: 0] pb_dma_to_descriptor_memory_s1_nativeaddress;
  output           pb_dma_to_descriptor_memory_s1_read;
  output  [ 31: 0] pb_dma_to_descriptor_memory_s1_readdata_from_sa;
  output           pb_dma_to_descriptor_memory_s1_reset_n;
  output           pb_dma_to_descriptor_memory_s1_waitrequest_from_sa;
  output           pb_dma_to_descriptor_memory_s1_write;
  output  [ 31: 0] pb_dma_to_descriptor_memory_s1_writedata;
  output           sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1;
  output           sgdma_rx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1;
  output           sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1;
  output           sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register;
  output           sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1;
  output           sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1;
  output           sgdma_rx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1;
  output           sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1;
  output           sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1;
  output           sgdma_tx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1;
  output           sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1;
  output           sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register;
  output           sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1;
  output           sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1;
  output           sgdma_tx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1;
  output           sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1;
  input            clk;
  input            pb_dma_to_descriptor_memory_s1_endofpacket;
  input   [ 31: 0] pb_dma_to_descriptor_memory_s1_readdata;
  input            pb_dma_to_descriptor_memory_s1_readdatavalid;
  input            pb_dma_to_descriptor_memory_s1_waitrequest;
  input            reset_n;
  input   [ 31: 0] sgdma_rx_descriptor_read_address_to_slave;
  input            sgdma_rx_descriptor_read_latency_counter;
  input            sgdma_rx_descriptor_read_read;
  input   [ 31: 0] sgdma_rx_descriptor_write_address_to_slave;
  input            sgdma_rx_descriptor_write_write;
  input   [ 31: 0] sgdma_rx_descriptor_write_writedata;
  input   [ 31: 0] sgdma_tx_descriptor_read_address_to_slave;
  input            sgdma_tx_descriptor_read_latency_counter;
  input            sgdma_tx_descriptor_read_read;
  input   [ 31: 0] sgdma_tx_descriptor_write_address_to_slave;
  input            sgdma_tx_descriptor_write_write;
  input   [ 31: 0] sgdma_tx_descriptor_write_writedata;

  reg              d1_pb_dma_to_descriptor_memory_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_pb_dma_to_descriptor_memory_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_sgdma_rx_descriptor_read_granted_slave_pb_dma_to_descriptor_memory_s1;
  reg              last_cycle_sgdma_rx_descriptor_write_granted_slave_pb_dma_to_descriptor_memory_s1;
  reg              last_cycle_sgdma_tx_descriptor_read_granted_slave_pb_dma_to_descriptor_memory_s1;
  reg              last_cycle_sgdma_tx_descriptor_write_granted_slave_pb_dma_to_descriptor_memory_s1;
  wire    [ 11: 0] pb_dma_to_descriptor_memory_s1_address;
  wire             pb_dma_to_descriptor_memory_s1_allgrants;
  wire             pb_dma_to_descriptor_memory_s1_allow_new_arb_cycle;
  wire             pb_dma_to_descriptor_memory_s1_any_bursting_master_saved_grant;
  wire             pb_dma_to_descriptor_memory_s1_any_continuerequest;
  reg     [  3: 0] pb_dma_to_descriptor_memory_s1_arb_addend;
  wire             pb_dma_to_descriptor_memory_s1_arb_counter_enable;
  reg     [  3: 0] pb_dma_to_descriptor_memory_s1_arb_share_counter;
  wire    [  3: 0] pb_dma_to_descriptor_memory_s1_arb_share_counter_next_value;
  wire    [  3: 0] pb_dma_to_descriptor_memory_s1_arb_share_set_values;
  wire    [  3: 0] pb_dma_to_descriptor_memory_s1_arb_winner;
  wire             pb_dma_to_descriptor_memory_s1_arbiterlock;
  wire             pb_dma_to_descriptor_memory_s1_arbiterlock2;
  wire             pb_dma_to_descriptor_memory_s1_arbitration_holdoff_internal;
  wire             pb_dma_to_descriptor_memory_s1_beginbursttransfer_internal;
  wire             pb_dma_to_descriptor_memory_s1_begins_xfer;
  wire             pb_dma_to_descriptor_memory_s1_burstcount;
  wire    [  3: 0] pb_dma_to_descriptor_memory_s1_byteenable;
  wire             pb_dma_to_descriptor_memory_s1_chipselect;
  wire    [  7: 0] pb_dma_to_descriptor_memory_s1_chosen_master_double_vector;
  wire    [  3: 0] pb_dma_to_descriptor_memory_s1_chosen_master_rot_left;
  wire             pb_dma_to_descriptor_memory_s1_debugaccess;
  wire             pb_dma_to_descriptor_memory_s1_end_xfer;
  wire             pb_dma_to_descriptor_memory_s1_endofpacket_from_sa;
  wire             pb_dma_to_descriptor_memory_s1_firsttransfer;
  wire    [  3: 0] pb_dma_to_descriptor_memory_s1_grant_vector;
  wire             pb_dma_to_descriptor_memory_s1_in_a_read_cycle;
  wire             pb_dma_to_descriptor_memory_s1_in_a_write_cycle;
  wire    [  3: 0] pb_dma_to_descriptor_memory_s1_master_qreq_vector;
  wire             pb_dma_to_descriptor_memory_s1_move_on_to_next_transaction;
  wire    [ 11: 0] pb_dma_to_descriptor_memory_s1_nativeaddress;
  wire             pb_dma_to_descriptor_memory_s1_non_bursting_master_requests;
  wire             pb_dma_to_descriptor_memory_s1_read;
  wire    [ 31: 0] pb_dma_to_descriptor_memory_s1_readdata_from_sa;
  wire             pb_dma_to_descriptor_memory_s1_readdatavalid_from_sa;
  reg              pb_dma_to_descriptor_memory_s1_reg_firsttransfer;
  wire             pb_dma_to_descriptor_memory_s1_reset_n;
  reg     [  3: 0] pb_dma_to_descriptor_memory_s1_saved_chosen_master_vector;
  reg              pb_dma_to_descriptor_memory_s1_slavearbiterlockenable;
  wire             pb_dma_to_descriptor_memory_s1_slavearbiterlockenable2;
  wire             pb_dma_to_descriptor_memory_s1_unreg_firsttransfer;
  wire             pb_dma_to_descriptor_memory_s1_waitrequest_from_sa;
  wire             pb_dma_to_descriptor_memory_s1_waits_for_read;
  wire             pb_dma_to_descriptor_memory_s1_waits_for_write;
  wire             pb_dma_to_descriptor_memory_s1_write;
  wire    [ 31: 0] pb_dma_to_descriptor_memory_s1_writedata;
  wire             sgdma_rx_descriptor_read_arbiterlock;
  wire             sgdma_rx_descriptor_read_arbiterlock2;
  wire             sgdma_rx_descriptor_read_continuerequest;
  wire             sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_rdv_fifo_empty_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_rdv_fifo_output_from_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register;
  wire             sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_saved_grant_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_arbiterlock;
  wire             sgdma_rx_descriptor_write_arbiterlock2;
  wire             sgdma_rx_descriptor_write_continuerequest;
  wire             sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_saved_grant_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_arbiterlock;
  wire             sgdma_tx_descriptor_read_arbiterlock2;
  wire             sgdma_tx_descriptor_read_continuerequest;
  wire             sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_rdv_fifo_empty_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_rdv_fifo_output_from_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register;
  wire             sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_saved_grant_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_arbiterlock;
  wire             sgdma_tx_descriptor_write_arbiterlock2;
  wire             sgdma_tx_descriptor_write_continuerequest;
  wire             sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_saved_grant_pb_dma_to_descriptor_memory_s1;
  wire    [ 31: 0] shifted_address_to_pb_dma_to_descriptor_memory_s1_from_sgdma_rx_descriptor_read;
  wire    [ 31: 0] shifted_address_to_pb_dma_to_descriptor_memory_s1_from_sgdma_rx_descriptor_write;
  wire    [ 31: 0] shifted_address_to_pb_dma_to_descriptor_memory_s1_from_sgdma_tx_descriptor_read;
  wire    [ 31: 0] shifted_address_to_pb_dma_to_descriptor_memory_s1_from_sgdma_tx_descriptor_write;
  wire             wait_for_pb_dma_to_descriptor_memory_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~pb_dma_to_descriptor_memory_s1_end_xfer;
    end


  assign pb_dma_to_descriptor_memory_s1_begins_xfer = ~d1_reasons_to_wait & ((sgdma_rx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1 | sgdma_rx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1 | sgdma_tx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1 | sgdma_tx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1));
  //assign pb_dma_to_descriptor_memory_s1_readdata_from_sa = pb_dma_to_descriptor_memory_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_readdata_from_sa = pb_dma_to_descriptor_memory_s1_readdata;

  assign sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1 = (({sgdma_rx_descriptor_read_address_to_slave[31 : 14] , 14'b0} == 32'h8000000) & (sgdma_rx_descriptor_read_read)) & sgdma_rx_descriptor_read_read;
  //assign pb_dma_to_descriptor_memory_s1_waitrequest_from_sa = pb_dma_to_descriptor_memory_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_waitrequest_from_sa = pb_dma_to_descriptor_memory_s1_waitrequest;

  //assign pb_dma_to_descriptor_memory_s1_readdatavalid_from_sa = pb_dma_to_descriptor_memory_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_readdatavalid_from_sa = pb_dma_to_descriptor_memory_s1_readdatavalid;

  //pb_dma_to_descriptor_memory_s1_arb_share_counter set values, which is an e_mux
  assign pb_dma_to_descriptor_memory_s1_arb_share_set_values = (sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1)? 8 :
    1;

  //pb_dma_to_descriptor_memory_s1_non_bursting_master_requests mux, which is an e_mux
  assign pb_dma_to_descriptor_memory_s1_non_bursting_master_requests = sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1 |
    sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1;

  //pb_dma_to_descriptor_memory_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign pb_dma_to_descriptor_memory_s1_any_bursting_master_saved_grant = 0;

  //pb_dma_to_descriptor_memory_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_arb_share_counter_next_value = pb_dma_to_descriptor_memory_s1_firsttransfer ? (pb_dma_to_descriptor_memory_s1_arb_share_set_values - 1) : |pb_dma_to_descriptor_memory_s1_arb_share_counter ? (pb_dma_to_descriptor_memory_s1_arb_share_counter - 1) : 0;

  //pb_dma_to_descriptor_memory_s1_allgrants all slave grants, which is an e_mux
  assign pb_dma_to_descriptor_memory_s1_allgrants = (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector) |
    (|pb_dma_to_descriptor_memory_s1_grant_vector);

  //pb_dma_to_descriptor_memory_s1_end_xfer assignment, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_end_xfer = ~(pb_dma_to_descriptor_memory_s1_waits_for_read | pb_dma_to_descriptor_memory_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_pb_dma_to_descriptor_memory_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_pb_dma_to_descriptor_memory_s1 = pb_dma_to_descriptor_memory_s1_end_xfer & (~pb_dma_to_descriptor_memory_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //pb_dma_to_descriptor_memory_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_pb_dma_to_descriptor_memory_s1 & pb_dma_to_descriptor_memory_s1_allgrants) | (end_xfer_arb_share_counter_term_pb_dma_to_descriptor_memory_s1 & ~pb_dma_to_descriptor_memory_s1_non_bursting_master_requests);

  //pb_dma_to_descriptor_memory_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_descriptor_memory_s1_arb_share_counter <= 0;
      else if (pb_dma_to_descriptor_memory_s1_arb_counter_enable)
          pb_dma_to_descriptor_memory_s1_arb_share_counter <= pb_dma_to_descriptor_memory_s1_arb_share_counter_next_value;
    end


  //pb_dma_to_descriptor_memory_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_descriptor_memory_s1_slavearbiterlockenable <= 0;
      else if ((|pb_dma_to_descriptor_memory_s1_master_qreq_vector & end_xfer_arb_share_counter_term_pb_dma_to_descriptor_memory_s1) | (end_xfer_arb_share_counter_term_pb_dma_to_descriptor_memory_s1 & ~pb_dma_to_descriptor_memory_s1_non_bursting_master_requests))
          pb_dma_to_descriptor_memory_s1_slavearbiterlockenable <= |pb_dma_to_descriptor_memory_s1_arb_share_counter_next_value;
    end


  //sgdma_rx/descriptor_read pb_dma_to_descriptor_memory/s1 arbiterlock, which is an e_assign
  assign sgdma_rx_descriptor_read_arbiterlock = pb_dma_to_descriptor_memory_s1_slavearbiterlockenable & sgdma_rx_descriptor_read_continuerequest;

  //pb_dma_to_descriptor_memory_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_slavearbiterlockenable2 = |pb_dma_to_descriptor_memory_s1_arb_share_counter_next_value;

  //sgdma_rx/descriptor_read pb_dma_to_descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign sgdma_rx_descriptor_read_arbiterlock2 = pb_dma_to_descriptor_memory_s1_slavearbiterlockenable2 & sgdma_rx_descriptor_read_continuerequest;

  //sgdma_rx/descriptor_write pb_dma_to_descriptor_memory/s1 arbiterlock, which is an e_assign
  assign sgdma_rx_descriptor_write_arbiterlock = pb_dma_to_descriptor_memory_s1_slavearbiterlockenable & sgdma_rx_descriptor_write_continuerequest;

  //sgdma_rx/descriptor_write pb_dma_to_descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign sgdma_rx_descriptor_write_arbiterlock2 = pb_dma_to_descriptor_memory_s1_slavearbiterlockenable2 & sgdma_rx_descriptor_write_continuerequest;

  //sgdma_rx/descriptor_write granted pb_dma_to_descriptor_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_rx_descriptor_write_granted_slave_pb_dma_to_descriptor_memory_s1 <= 0;
      else 
        last_cycle_sgdma_rx_descriptor_write_granted_slave_pb_dma_to_descriptor_memory_s1 <= sgdma_rx_descriptor_write_saved_grant_pb_dma_to_descriptor_memory_s1 ? 1 : (pb_dma_to_descriptor_memory_s1_arbitration_holdoff_internal | ~sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1) ? 0 : last_cycle_sgdma_rx_descriptor_write_granted_slave_pb_dma_to_descriptor_memory_s1;
    end


  //sgdma_rx_descriptor_write_continuerequest continued request, which is an e_mux
  assign sgdma_rx_descriptor_write_continuerequest = (last_cycle_sgdma_rx_descriptor_write_granted_slave_pb_dma_to_descriptor_memory_s1 & sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_write_granted_slave_pb_dma_to_descriptor_memory_s1 & sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_write_granted_slave_pb_dma_to_descriptor_memory_s1 & sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1);

  //pb_dma_to_descriptor_memory_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign pb_dma_to_descriptor_memory_s1_any_continuerequest = sgdma_rx_descriptor_write_continuerequest |
    sgdma_tx_descriptor_read_continuerequest |
    sgdma_tx_descriptor_write_continuerequest |
    sgdma_rx_descriptor_read_continuerequest |
    sgdma_tx_descriptor_read_continuerequest |
    sgdma_tx_descriptor_write_continuerequest |
    sgdma_rx_descriptor_read_continuerequest |
    sgdma_rx_descriptor_write_continuerequest |
    sgdma_tx_descriptor_write_continuerequest |
    sgdma_rx_descriptor_read_continuerequest |
    sgdma_rx_descriptor_write_continuerequest |
    sgdma_tx_descriptor_read_continuerequest;

  //sgdma_tx/descriptor_read pb_dma_to_descriptor_memory/s1 arbiterlock, which is an e_assign
  assign sgdma_tx_descriptor_read_arbiterlock = pb_dma_to_descriptor_memory_s1_slavearbiterlockenable & sgdma_tx_descriptor_read_continuerequest;

  //sgdma_tx/descriptor_read pb_dma_to_descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign sgdma_tx_descriptor_read_arbiterlock2 = pb_dma_to_descriptor_memory_s1_slavearbiterlockenable2 & sgdma_tx_descriptor_read_continuerequest;

  //sgdma_tx/descriptor_read granted pb_dma_to_descriptor_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_tx_descriptor_read_granted_slave_pb_dma_to_descriptor_memory_s1 <= 0;
      else 
        last_cycle_sgdma_tx_descriptor_read_granted_slave_pb_dma_to_descriptor_memory_s1 <= sgdma_tx_descriptor_read_saved_grant_pb_dma_to_descriptor_memory_s1 ? 1 : (pb_dma_to_descriptor_memory_s1_arbitration_holdoff_internal | ~sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1) ? 0 : last_cycle_sgdma_tx_descriptor_read_granted_slave_pb_dma_to_descriptor_memory_s1;
    end


  //sgdma_tx_descriptor_read_continuerequest continued request, which is an e_mux
  assign sgdma_tx_descriptor_read_continuerequest = (last_cycle_sgdma_tx_descriptor_read_granted_slave_pb_dma_to_descriptor_memory_s1 & sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_read_granted_slave_pb_dma_to_descriptor_memory_s1 & sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_read_granted_slave_pb_dma_to_descriptor_memory_s1 & sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1);

  //sgdma_tx/descriptor_write pb_dma_to_descriptor_memory/s1 arbiterlock, which is an e_assign
  assign sgdma_tx_descriptor_write_arbiterlock = pb_dma_to_descriptor_memory_s1_slavearbiterlockenable & sgdma_tx_descriptor_write_continuerequest;

  //sgdma_tx/descriptor_write pb_dma_to_descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign sgdma_tx_descriptor_write_arbiterlock2 = pb_dma_to_descriptor_memory_s1_slavearbiterlockenable2 & sgdma_tx_descriptor_write_continuerequest;

  //sgdma_tx/descriptor_write granted pb_dma_to_descriptor_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_tx_descriptor_write_granted_slave_pb_dma_to_descriptor_memory_s1 <= 0;
      else 
        last_cycle_sgdma_tx_descriptor_write_granted_slave_pb_dma_to_descriptor_memory_s1 <= sgdma_tx_descriptor_write_saved_grant_pb_dma_to_descriptor_memory_s1 ? 1 : (pb_dma_to_descriptor_memory_s1_arbitration_holdoff_internal | ~sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1) ? 0 : last_cycle_sgdma_tx_descriptor_write_granted_slave_pb_dma_to_descriptor_memory_s1;
    end


  //sgdma_tx_descriptor_write_continuerequest continued request, which is an e_mux
  assign sgdma_tx_descriptor_write_continuerequest = (last_cycle_sgdma_tx_descriptor_write_granted_slave_pb_dma_to_descriptor_memory_s1 & sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_write_granted_slave_pb_dma_to_descriptor_memory_s1 & sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_write_granted_slave_pb_dma_to_descriptor_memory_s1 & sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1);

  assign sgdma_rx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1 = sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1 & ~((sgdma_rx_descriptor_read_read & ((sgdma_rx_descriptor_read_latency_counter != 0) | (1 < sgdma_rx_descriptor_read_latency_counter))) | sgdma_rx_descriptor_write_arbiterlock | sgdma_tx_descriptor_read_arbiterlock | sgdma_tx_descriptor_write_arbiterlock);
  //unique name for pb_dma_to_descriptor_memory_s1_move_on_to_next_transaction, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_move_on_to_next_transaction = pb_dma_to_descriptor_memory_s1_readdatavalid_from_sa;

  //rdv_fifo_for_sgdma_rx_descriptor_read_to_pb_dma_to_descriptor_memory_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_sgdma_rx_descriptor_read_to_pb_dma_to_descriptor_memory_s1_module rdv_fifo_for_sgdma_rx_descriptor_read_to_pb_dma_to_descriptor_memory_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1),
      .data_out             (sgdma_rx_descriptor_read_rdv_fifo_output_from_pb_dma_to_descriptor_memory_s1),
      .empty                (),
      .fifo_contains_ones_n (sgdma_rx_descriptor_read_rdv_fifo_empty_pb_dma_to_descriptor_memory_s1),
      .full                 (),
      .read                 (pb_dma_to_descriptor_memory_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~pb_dma_to_descriptor_memory_s1_waits_for_read)
    );

  assign sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register = ~sgdma_rx_descriptor_read_rdv_fifo_empty_pb_dma_to_descriptor_memory_s1;
  //local readdatavalid sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1, which is an e_mux
  assign sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1 = (pb_dma_to_descriptor_memory_s1_readdatavalid_from_sa & sgdma_rx_descriptor_read_rdv_fifo_output_from_pb_dma_to_descriptor_memory_s1) & ~ sgdma_rx_descriptor_read_rdv_fifo_empty_pb_dma_to_descriptor_memory_s1;

  //assign pb_dma_to_descriptor_memory_s1_endofpacket_from_sa = pb_dma_to_descriptor_memory_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_endofpacket_from_sa = pb_dma_to_descriptor_memory_s1_endofpacket;

  assign sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1 = (({sgdma_rx_descriptor_write_address_to_slave[31 : 14] , 14'b0} == 32'h8000000) & (sgdma_rx_descriptor_write_write)) & sgdma_rx_descriptor_write_write;
  //sgdma_rx/descriptor_read granted pb_dma_to_descriptor_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_rx_descriptor_read_granted_slave_pb_dma_to_descriptor_memory_s1 <= 0;
      else 
        last_cycle_sgdma_rx_descriptor_read_granted_slave_pb_dma_to_descriptor_memory_s1 <= sgdma_rx_descriptor_read_saved_grant_pb_dma_to_descriptor_memory_s1 ? 1 : (pb_dma_to_descriptor_memory_s1_arbitration_holdoff_internal | ~sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1) ? 0 : last_cycle_sgdma_rx_descriptor_read_granted_slave_pb_dma_to_descriptor_memory_s1;
    end


  //sgdma_rx_descriptor_read_continuerequest continued request, which is an e_mux
  assign sgdma_rx_descriptor_read_continuerequest = (last_cycle_sgdma_rx_descriptor_read_granted_slave_pb_dma_to_descriptor_memory_s1 & sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_read_granted_slave_pb_dma_to_descriptor_memory_s1 & sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_read_granted_slave_pb_dma_to_descriptor_memory_s1 & sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1);

  assign sgdma_rx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1 = sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1 & ~(sgdma_rx_descriptor_read_arbiterlock | sgdma_tx_descriptor_read_arbiterlock | sgdma_tx_descriptor_write_arbiterlock);
  //pb_dma_to_descriptor_memory_s1_writedata mux, which is an e_mux
  assign pb_dma_to_descriptor_memory_s1_writedata = (sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1)? sgdma_rx_descriptor_write_writedata :
    sgdma_tx_descriptor_write_writedata;

  assign sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1 = (({sgdma_tx_descriptor_read_address_to_slave[31 : 14] , 14'b0} == 32'h8000000) & (sgdma_tx_descriptor_read_read)) & sgdma_tx_descriptor_read_read;
  assign sgdma_tx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1 = sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1 & ~((sgdma_tx_descriptor_read_read & ((sgdma_tx_descriptor_read_latency_counter != 0) | (1 < sgdma_tx_descriptor_read_latency_counter))) | sgdma_rx_descriptor_read_arbiterlock | sgdma_rx_descriptor_write_arbiterlock | sgdma_tx_descriptor_write_arbiterlock);
  //rdv_fifo_for_sgdma_tx_descriptor_read_to_pb_dma_to_descriptor_memory_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_sgdma_tx_descriptor_read_to_pb_dma_to_descriptor_memory_s1_module rdv_fifo_for_sgdma_tx_descriptor_read_to_pb_dma_to_descriptor_memory_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1),
      .data_out             (sgdma_tx_descriptor_read_rdv_fifo_output_from_pb_dma_to_descriptor_memory_s1),
      .empty                (),
      .fifo_contains_ones_n (sgdma_tx_descriptor_read_rdv_fifo_empty_pb_dma_to_descriptor_memory_s1),
      .full                 (),
      .read                 (pb_dma_to_descriptor_memory_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~pb_dma_to_descriptor_memory_s1_waits_for_read)
    );

  assign sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register = ~sgdma_tx_descriptor_read_rdv_fifo_empty_pb_dma_to_descriptor_memory_s1;
  //local readdatavalid sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1, which is an e_mux
  assign sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1 = (pb_dma_to_descriptor_memory_s1_readdatavalid_from_sa & sgdma_tx_descriptor_read_rdv_fifo_output_from_pb_dma_to_descriptor_memory_s1) & ~ sgdma_tx_descriptor_read_rdv_fifo_empty_pb_dma_to_descriptor_memory_s1;

  assign sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1 = (({sgdma_tx_descriptor_write_address_to_slave[31 : 14] , 14'b0} == 32'h8000000) & (sgdma_tx_descriptor_write_write)) & sgdma_tx_descriptor_write_write;
  assign sgdma_tx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1 = sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1 & ~(sgdma_rx_descriptor_read_arbiterlock | sgdma_rx_descriptor_write_arbiterlock | sgdma_tx_descriptor_read_arbiterlock);
  //allow new arb cycle for pb_dma_to_descriptor_memory/s1, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_allow_new_arb_cycle = ~sgdma_rx_descriptor_read_arbiterlock & ~sgdma_rx_descriptor_write_arbiterlock & ~sgdma_tx_descriptor_read_arbiterlock & ~sgdma_tx_descriptor_write_arbiterlock;

  //sgdma_tx/descriptor_write assignment into master qualified-requests vector for pb_dma_to_descriptor_memory/s1, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_master_qreq_vector[0] = sgdma_tx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1;

  //sgdma_tx/descriptor_write grant pb_dma_to_descriptor_memory/s1, which is an e_assign
  assign sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1 = pb_dma_to_descriptor_memory_s1_grant_vector[0];

  //sgdma_tx/descriptor_write saved-grant pb_dma_to_descriptor_memory/s1, which is an e_assign
  assign sgdma_tx_descriptor_write_saved_grant_pb_dma_to_descriptor_memory_s1 = pb_dma_to_descriptor_memory_s1_arb_winner[0] && sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1;

  //sgdma_tx/descriptor_read assignment into master qualified-requests vector for pb_dma_to_descriptor_memory/s1, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_master_qreq_vector[1] = sgdma_tx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1;

  //sgdma_tx/descriptor_read grant pb_dma_to_descriptor_memory/s1, which is an e_assign
  assign sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1 = pb_dma_to_descriptor_memory_s1_grant_vector[1];

  //sgdma_tx/descriptor_read saved-grant pb_dma_to_descriptor_memory/s1, which is an e_assign
  assign sgdma_tx_descriptor_read_saved_grant_pb_dma_to_descriptor_memory_s1 = pb_dma_to_descriptor_memory_s1_arb_winner[1] && sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1;

  //sgdma_rx/descriptor_write assignment into master qualified-requests vector for pb_dma_to_descriptor_memory/s1, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_master_qreq_vector[2] = sgdma_rx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1;

  //sgdma_rx/descriptor_write grant pb_dma_to_descriptor_memory/s1, which is an e_assign
  assign sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1 = pb_dma_to_descriptor_memory_s1_grant_vector[2];

  //sgdma_rx/descriptor_write saved-grant pb_dma_to_descriptor_memory/s1, which is an e_assign
  assign sgdma_rx_descriptor_write_saved_grant_pb_dma_to_descriptor_memory_s1 = pb_dma_to_descriptor_memory_s1_arb_winner[2] && sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1;

  //sgdma_rx/descriptor_read assignment into master qualified-requests vector for pb_dma_to_descriptor_memory/s1, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_master_qreq_vector[3] = sgdma_rx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1;

  //sgdma_rx/descriptor_read grant pb_dma_to_descriptor_memory/s1, which is an e_assign
  assign sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1 = pb_dma_to_descriptor_memory_s1_grant_vector[3];

  //sgdma_rx/descriptor_read saved-grant pb_dma_to_descriptor_memory/s1, which is an e_assign
  assign sgdma_rx_descriptor_read_saved_grant_pb_dma_to_descriptor_memory_s1 = pb_dma_to_descriptor_memory_s1_arb_winner[3] && sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1;

  //pb_dma_to_descriptor_memory/s1 chosen-master double-vector, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_chosen_master_double_vector = {pb_dma_to_descriptor_memory_s1_master_qreq_vector, pb_dma_to_descriptor_memory_s1_master_qreq_vector} & ({~pb_dma_to_descriptor_memory_s1_master_qreq_vector, ~pb_dma_to_descriptor_memory_s1_master_qreq_vector} + pb_dma_to_descriptor_memory_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign pb_dma_to_descriptor_memory_s1_arb_winner = (pb_dma_to_descriptor_memory_s1_allow_new_arb_cycle & | pb_dma_to_descriptor_memory_s1_grant_vector) ? pb_dma_to_descriptor_memory_s1_grant_vector : pb_dma_to_descriptor_memory_s1_saved_chosen_master_vector;

  //saved pb_dma_to_descriptor_memory_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_descriptor_memory_s1_saved_chosen_master_vector <= 0;
      else if (pb_dma_to_descriptor_memory_s1_allow_new_arb_cycle)
          pb_dma_to_descriptor_memory_s1_saved_chosen_master_vector <= |pb_dma_to_descriptor_memory_s1_grant_vector ? pb_dma_to_descriptor_memory_s1_grant_vector : pb_dma_to_descriptor_memory_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign pb_dma_to_descriptor_memory_s1_grant_vector = {(pb_dma_to_descriptor_memory_s1_chosen_master_double_vector[3] | pb_dma_to_descriptor_memory_s1_chosen_master_double_vector[7]),
    (pb_dma_to_descriptor_memory_s1_chosen_master_double_vector[2] | pb_dma_to_descriptor_memory_s1_chosen_master_double_vector[6]),
    (pb_dma_to_descriptor_memory_s1_chosen_master_double_vector[1] | pb_dma_to_descriptor_memory_s1_chosen_master_double_vector[5]),
    (pb_dma_to_descriptor_memory_s1_chosen_master_double_vector[0] | pb_dma_to_descriptor_memory_s1_chosen_master_double_vector[4])};

  //pb_dma_to_descriptor_memory/s1 chosen master rotated left, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_chosen_master_rot_left = (pb_dma_to_descriptor_memory_s1_arb_winner << 1) ? (pb_dma_to_descriptor_memory_s1_arb_winner << 1) : 1;

  //pb_dma_to_descriptor_memory/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_descriptor_memory_s1_arb_addend <= 1;
      else if (|pb_dma_to_descriptor_memory_s1_grant_vector)
          pb_dma_to_descriptor_memory_s1_arb_addend <= pb_dma_to_descriptor_memory_s1_end_xfer? pb_dma_to_descriptor_memory_s1_chosen_master_rot_left : pb_dma_to_descriptor_memory_s1_grant_vector;
    end


  //pb_dma_to_descriptor_memory_s1_reset_n assignment, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_reset_n = reset_n;

  assign pb_dma_to_descriptor_memory_s1_chipselect = sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1 | sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1 | sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1 | sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1;
  //pb_dma_to_descriptor_memory_s1_firsttransfer first transaction, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_firsttransfer = pb_dma_to_descriptor_memory_s1_begins_xfer ? pb_dma_to_descriptor_memory_s1_unreg_firsttransfer : pb_dma_to_descriptor_memory_s1_reg_firsttransfer;

  //pb_dma_to_descriptor_memory_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_unreg_firsttransfer = ~(pb_dma_to_descriptor_memory_s1_slavearbiterlockenable & pb_dma_to_descriptor_memory_s1_any_continuerequest);

  //pb_dma_to_descriptor_memory_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_descriptor_memory_s1_reg_firsttransfer <= 1'b1;
      else if (pb_dma_to_descriptor_memory_s1_begins_xfer)
          pb_dma_to_descriptor_memory_s1_reg_firsttransfer <= pb_dma_to_descriptor_memory_s1_unreg_firsttransfer;
    end


  //pb_dma_to_descriptor_memory_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_beginbursttransfer_internal = pb_dma_to_descriptor_memory_s1_begins_xfer;

  //pb_dma_to_descriptor_memory_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_arbitration_holdoff_internal = pb_dma_to_descriptor_memory_s1_begins_xfer & pb_dma_to_descriptor_memory_s1_firsttransfer;

  //pb_dma_to_descriptor_memory_s1_read assignment, which is an e_mux
  assign pb_dma_to_descriptor_memory_s1_read = (sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1 & sgdma_rx_descriptor_read_read) | (sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1 & sgdma_tx_descriptor_read_read);

  //pb_dma_to_descriptor_memory_s1_write assignment, which is an e_mux
  assign pb_dma_to_descriptor_memory_s1_write = (sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1 & sgdma_rx_descriptor_write_write) | (sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1 & sgdma_tx_descriptor_write_write);

  assign shifted_address_to_pb_dma_to_descriptor_memory_s1_from_sgdma_rx_descriptor_read = sgdma_rx_descriptor_read_address_to_slave;
  //pb_dma_to_descriptor_memory_s1_address mux, which is an e_mux
  assign pb_dma_to_descriptor_memory_s1_address = (sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1)? (shifted_address_to_pb_dma_to_descriptor_memory_s1_from_sgdma_rx_descriptor_read >> 2) :
    (sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1)? (shifted_address_to_pb_dma_to_descriptor_memory_s1_from_sgdma_rx_descriptor_write >> 2) :
    (sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1)? (shifted_address_to_pb_dma_to_descriptor_memory_s1_from_sgdma_tx_descriptor_read >> 2) :
    (shifted_address_to_pb_dma_to_descriptor_memory_s1_from_sgdma_tx_descriptor_write >> 2);

  assign shifted_address_to_pb_dma_to_descriptor_memory_s1_from_sgdma_rx_descriptor_write = sgdma_rx_descriptor_write_address_to_slave;
  assign shifted_address_to_pb_dma_to_descriptor_memory_s1_from_sgdma_tx_descriptor_read = sgdma_tx_descriptor_read_address_to_slave;
  assign shifted_address_to_pb_dma_to_descriptor_memory_s1_from_sgdma_tx_descriptor_write = sgdma_tx_descriptor_write_address_to_slave;
  //slaveid pb_dma_to_descriptor_memory_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign pb_dma_to_descriptor_memory_s1_nativeaddress = (sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1)? (sgdma_rx_descriptor_read_address_to_slave >> 2) :
    (sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1)? (sgdma_rx_descriptor_write_address_to_slave >> 2) :
    (sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1)? (sgdma_tx_descriptor_read_address_to_slave >> 2) :
    (sgdma_tx_descriptor_write_address_to_slave >> 2);

  //d1_pb_dma_to_descriptor_memory_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_pb_dma_to_descriptor_memory_s1_end_xfer <= 1;
      else 
        d1_pb_dma_to_descriptor_memory_s1_end_xfer <= pb_dma_to_descriptor_memory_s1_end_xfer;
    end


  //pb_dma_to_descriptor_memory_s1_waits_for_read in a cycle, which is an e_mux
  assign pb_dma_to_descriptor_memory_s1_waits_for_read = pb_dma_to_descriptor_memory_s1_in_a_read_cycle & pb_dma_to_descriptor_memory_s1_waitrequest_from_sa;

  //pb_dma_to_descriptor_memory_s1_in_a_read_cycle assignment, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_in_a_read_cycle = (sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1 & sgdma_rx_descriptor_read_read) | (sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1 & sgdma_tx_descriptor_read_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = pb_dma_to_descriptor_memory_s1_in_a_read_cycle;

  //pb_dma_to_descriptor_memory_s1_waits_for_write in a cycle, which is an e_mux
  assign pb_dma_to_descriptor_memory_s1_waits_for_write = pb_dma_to_descriptor_memory_s1_in_a_write_cycle & pb_dma_to_descriptor_memory_s1_waitrequest_from_sa;

  //pb_dma_to_descriptor_memory_s1_in_a_write_cycle assignment, which is an e_assign
  assign pb_dma_to_descriptor_memory_s1_in_a_write_cycle = (sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1 & sgdma_rx_descriptor_write_write) | (sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1 & sgdma_tx_descriptor_write_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = pb_dma_to_descriptor_memory_s1_in_a_write_cycle;

  assign wait_for_pb_dma_to_descriptor_memory_s1_counter = 0;
  //pb_dma_to_descriptor_memory_s1_byteenable byte enable port mux, which is an e_mux
  assign pb_dma_to_descriptor_memory_s1_byteenable = (sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1)? {4 {1'b1}} :
    (sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1)? {4 {1'b1}} :
    -1;

  //burstcount mux, which is an e_mux
  assign pb_dma_to_descriptor_memory_s1_burstcount = 1;

  //pb_dma_to_descriptor_memory/s1 arbiterlock assigned from _handle_arbiterlock, which is an e_mux
  assign pb_dma_to_descriptor_memory_s1_arbiterlock = (sgdma_rx_descriptor_read_arbiterlock)? sgdma_rx_descriptor_read_arbiterlock :
    (sgdma_rx_descriptor_write_arbiterlock)? sgdma_rx_descriptor_write_arbiterlock :
    (sgdma_tx_descriptor_read_arbiterlock)? sgdma_tx_descriptor_read_arbiterlock :
    sgdma_tx_descriptor_write_arbiterlock;

  //pb_dma_to_descriptor_memory/s1 arbiterlock2 assigned from _handle_arbiterlock2, which is an e_mux
  assign pb_dma_to_descriptor_memory_s1_arbiterlock2 = (sgdma_rx_descriptor_read_arbiterlock2)? sgdma_rx_descriptor_read_arbiterlock2 :
    (sgdma_rx_descriptor_write_arbiterlock2)? sgdma_rx_descriptor_write_arbiterlock2 :
    (sgdma_tx_descriptor_read_arbiterlock2)? sgdma_tx_descriptor_read_arbiterlock2 :
    sgdma_tx_descriptor_write_arbiterlock2;

  //debugaccess mux, which is an e_mux
  assign pb_dma_to_descriptor_memory_s1_debugaccess = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pb_dma_to_descriptor_memory/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1 + sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1 + sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1 + sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (sgdma_rx_descriptor_read_saved_grant_pb_dma_to_descriptor_memory_s1 + sgdma_rx_descriptor_write_saved_grant_pb_dma_to_descriptor_memory_s1 + sgdma_tx_descriptor_read_saved_grant_pb_dma_to_descriptor_memory_s1 + sgdma_tx_descriptor_write_saved_grant_pb_dma_to_descriptor_memory_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pb_dma_to_descriptor_memory_m1_arbitrator (
                                                   // inputs:
                                                    clk,
                                                    d1_descriptor_memory_s1_end_xfer,
                                                    descriptor_memory_s1_readdata_from_sa,
                                                    pb_dma_to_descriptor_memory_m1_address,
                                                    pb_dma_to_descriptor_memory_m1_burstcount,
                                                    pb_dma_to_descriptor_memory_m1_byteenable,
                                                    pb_dma_to_descriptor_memory_m1_chipselect,
                                                    pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1,
                                                    pb_dma_to_descriptor_memory_m1_qualified_request_descriptor_memory_s1,
                                                    pb_dma_to_descriptor_memory_m1_read,
                                                    pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1,
                                                    pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1,
                                                    pb_dma_to_descriptor_memory_m1_write,
                                                    pb_dma_to_descriptor_memory_m1_writedata,
                                                    reset_n,

                                                   // outputs:
                                                    pb_dma_to_descriptor_memory_m1_address_to_slave,
                                                    pb_dma_to_descriptor_memory_m1_latency_counter,
                                                    pb_dma_to_descriptor_memory_m1_readdata,
                                                    pb_dma_to_descriptor_memory_m1_readdatavalid,
                                                    pb_dma_to_descriptor_memory_m1_waitrequest
                                                 )
;

  output  [ 13: 0] pb_dma_to_descriptor_memory_m1_address_to_slave;
  output           pb_dma_to_descriptor_memory_m1_latency_counter;
  output  [ 31: 0] pb_dma_to_descriptor_memory_m1_readdata;
  output           pb_dma_to_descriptor_memory_m1_readdatavalid;
  output           pb_dma_to_descriptor_memory_m1_waitrequest;
  input            clk;
  input            d1_descriptor_memory_s1_end_xfer;
  input   [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  input   [ 13: 0] pb_dma_to_descriptor_memory_m1_address;
  input            pb_dma_to_descriptor_memory_m1_burstcount;
  input   [  3: 0] pb_dma_to_descriptor_memory_m1_byteenable;
  input            pb_dma_to_descriptor_memory_m1_chipselect;
  input            pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1;
  input            pb_dma_to_descriptor_memory_m1_qualified_request_descriptor_memory_s1;
  input            pb_dma_to_descriptor_memory_m1_read;
  input            pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1;
  input            pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1;
  input            pb_dma_to_descriptor_memory_m1_write;
  input   [ 31: 0] pb_dma_to_descriptor_memory_m1_writedata;
  input            reset_n;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_pb_dma_to_descriptor_memory_m1_latency_counter;
  reg     [ 13: 0] pb_dma_to_descriptor_memory_m1_address_last_time;
  wire    [ 13: 0] pb_dma_to_descriptor_memory_m1_address_to_slave;
  reg              pb_dma_to_descriptor_memory_m1_burstcount_last_time;
  reg     [  3: 0] pb_dma_to_descriptor_memory_m1_byteenable_last_time;
  reg              pb_dma_to_descriptor_memory_m1_chipselect_last_time;
  wire             pb_dma_to_descriptor_memory_m1_is_granted_some_slave;
  reg              pb_dma_to_descriptor_memory_m1_latency_counter;
  reg              pb_dma_to_descriptor_memory_m1_read_but_no_slave_selected;
  reg              pb_dma_to_descriptor_memory_m1_read_last_time;
  wire    [ 31: 0] pb_dma_to_descriptor_memory_m1_readdata;
  wire             pb_dma_to_descriptor_memory_m1_readdatavalid;
  wire             pb_dma_to_descriptor_memory_m1_run;
  wire             pb_dma_to_descriptor_memory_m1_waitrequest;
  reg              pb_dma_to_descriptor_memory_m1_write_last_time;
  reg     [ 31: 0] pb_dma_to_descriptor_memory_m1_writedata_last_time;
  wire             pre_flush_pb_dma_to_descriptor_memory_m1_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (pb_dma_to_descriptor_memory_m1_qualified_request_descriptor_memory_s1 | ~pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1) & (pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1 | ~pb_dma_to_descriptor_memory_m1_qualified_request_descriptor_memory_s1) & ((~pb_dma_to_descriptor_memory_m1_qualified_request_descriptor_memory_s1 | ~pb_dma_to_descriptor_memory_m1_chipselect | (1 & pb_dma_to_descriptor_memory_m1_chipselect))) & ((~pb_dma_to_descriptor_memory_m1_qualified_request_descriptor_memory_s1 | ~pb_dma_to_descriptor_memory_m1_chipselect | (1 & pb_dma_to_descriptor_memory_m1_chipselect)));

  //cascaded wait assignment, which is an e_assign
  assign pb_dma_to_descriptor_memory_m1_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign pb_dma_to_descriptor_memory_m1_address_to_slave = {1'b1,
    pb_dma_to_descriptor_memory_m1_address[12 : 0]};

  //pb_dma_to_descriptor_memory_m1_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_descriptor_memory_m1_read_but_no_slave_selected <= 0;
      else 
        pb_dma_to_descriptor_memory_m1_read_but_no_slave_selected <= (pb_dma_to_descriptor_memory_m1_read & pb_dma_to_descriptor_memory_m1_chipselect) & pb_dma_to_descriptor_memory_m1_run & ~pb_dma_to_descriptor_memory_m1_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign pb_dma_to_descriptor_memory_m1_is_granted_some_slave = pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_pb_dma_to_descriptor_memory_m1_readdatavalid = pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign pb_dma_to_descriptor_memory_m1_readdatavalid = pb_dma_to_descriptor_memory_m1_read_but_no_slave_selected |
    pre_flush_pb_dma_to_descriptor_memory_m1_readdatavalid;

  //pb_dma_to_descriptor_memory/m1 readdata mux, which is an e_mux
  assign pb_dma_to_descriptor_memory_m1_readdata = descriptor_memory_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign pb_dma_to_descriptor_memory_m1_waitrequest = ~pb_dma_to_descriptor_memory_m1_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_descriptor_memory_m1_latency_counter <= 0;
      else 
        pb_dma_to_descriptor_memory_m1_latency_counter <= p1_pb_dma_to_descriptor_memory_m1_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_pb_dma_to_descriptor_memory_m1_latency_counter = ((pb_dma_to_descriptor_memory_m1_run & (pb_dma_to_descriptor_memory_m1_read & pb_dma_to_descriptor_memory_m1_chipselect)))? latency_load_value :
    (pb_dma_to_descriptor_memory_m1_latency_counter)? pb_dma_to_descriptor_memory_m1_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {1 {pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1}} & 1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pb_dma_to_descriptor_memory_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_descriptor_memory_m1_address_last_time <= 0;
      else 
        pb_dma_to_descriptor_memory_m1_address_last_time <= pb_dma_to_descriptor_memory_m1_address;
    end


  //pb_dma_to_descriptor_memory/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= pb_dma_to_descriptor_memory_m1_waitrequest & pb_dma_to_descriptor_memory_m1_chipselect;
    end


  //pb_dma_to_descriptor_memory_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_dma_to_descriptor_memory_m1_address != pb_dma_to_descriptor_memory_m1_address_last_time))
        begin
          $write("%0d ns: pb_dma_to_descriptor_memory_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_dma_to_descriptor_memory_m1_chipselect check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_descriptor_memory_m1_chipselect_last_time <= 0;
      else 
        pb_dma_to_descriptor_memory_m1_chipselect_last_time <= pb_dma_to_descriptor_memory_m1_chipselect;
    end


  //pb_dma_to_descriptor_memory_m1_chipselect matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_dma_to_descriptor_memory_m1_chipselect != pb_dma_to_descriptor_memory_m1_chipselect_last_time))
        begin
          $write("%0d ns: pb_dma_to_descriptor_memory_m1_chipselect did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_dma_to_descriptor_memory_m1_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_descriptor_memory_m1_burstcount_last_time <= 0;
      else 
        pb_dma_to_descriptor_memory_m1_burstcount_last_time <= pb_dma_to_descriptor_memory_m1_burstcount;
    end


  //pb_dma_to_descriptor_memory_m1_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_dma_to_descriptor_memory_m1_burstcount != pb_dma_to_descriptor_memory_m1_burstcount_last_time))
        begin
          $write("%0d ns: pb_dma_to_descriptor_memory_m1_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_dma_to_descriptor_memory_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_descriptor_memory_m1_byteenable_last_time <= 0;
      else 
        pb_dma_to_descriptor_memory_m1_byteenable_last_time <= pb_dma_to_descriptor_memory_m1_byteenable;
    end


  //pb_dma_to_descriptor_memory_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_dma_to_descriptor_memory_m1_byteenable != pb_dma_to_descriptor_memory_m1_byteenable_last_time))
        begin
          $write("%0d ns: pb_dma_to_descriptor_memory_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_dma_to_descriptor_memory_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_descriptor_memory_m1_read_last_time <= 0;
      else 
        pb_dma_to_descriptor_memory_m1_read_last_time <= pb_dma_to_descriptor_memory_m1_read;
    end


  //pb_dma_to_descriptor_memory_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_dma_to_descriptor_memory_m1_read != pb_dma_to_descriptor_memory_m1_read_last_time))
        begin
          $write("%0d ns: pb_dma_to_descriptor_memory_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_dma_to_descriptor_memory_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_descriptor_memory_m1_write_last_time <= 0;
      else 
        pb_dma_to_descriptor_memory_m1_write_last_time <= pb_dma_to_descriptor_memory_m1_write;
    end


  //pb_dma_to_descriptor_memory_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_dma_to_descriptor_memory_m1_write != pb_dma_to_descriptor_memory_m1_write_last_time))
        begin
          $write("%0d ns: pb_dma_to_descriptor_memory_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //pb_dma_to_descriptor_memory_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_dma_to_descriptor_memory_m1_writedata_last_time <= 0;
      else 
        pb_dma_to_descriptor_memory_m1_writedata_last_time <= pb_dma_to_descriptor_memory_m1_writedata;
    end


  //pb_dma_to_descriptor_memory_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pb_dma_to_descriptor_memory_m1_writedata != pb_dma_to_descriptor_memory_m1_writedata_last_time) & (pb_dma_to_descriptor_memory_m1_write & pb_dma_to_descriptor_memory_m1_chipselect))
        begin
          $write("%0d ns: pb_dma_to_descriptor_memory_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pb_dma_to_descriptor_memory_bridge_arbitrator 
;



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_rx_csr_arbitrator (
                                 // inputs:
                                  clk,
                                  pb_cpu_to_io_m1_address_to_slave,
                                  pb_cpu_to_io_m1_burstcount,
                                  pb_cpu_to_io_m1_chipselect,
                                  pb_cpu_to_io_m1_latency_counter,
                                  pb_cpu_to_io_m1_read,
                                  pb_cpu_to_io_m1_write,
                                  pb_cpu_to_io_m1_writedata,
                                  reset_n,
                                  sgdma_rx_csr_irq,
                                  sgdma_rx_csr_readdata,

                                 // outputs:
                                  d1_sgdma_rx_csr_end_xfer,
                                  pb_cpu_to_io_m1_granted_sgdma_rx_csr,
                                  pb_cpu_to_io_m1_qualified_request_sgdma_rx_csr,
                                  pb_cpu_to_io_m1_read_data_valid_sgdma_rx_csr,
                                  pb_cpu_to_io_m1_requests_sgdma_rx_csr,
                                  sgdma_rx_csr_address,
                                  sgdma_rx_csr_chipselect,
                                  sgdma_rx_csr_irq_from_sa,
                                  sgdma_rx_csr_read,
                                  sgdma_rx_csr_readdata_from_sa,
                                  sgdma_rx_csr_reset_n,
                                  sgdma_rx_csr_write,
                                  sgdma_rx_csr_writedata
                               )
;

  output           d1_sgdma_rx_csr_end_xfer;
  output           pb_cpu_to_io_m1_granted_sgdma_rx_csr;
  output           pb_cpu_to_io_m1_qualified_request_sgdma_rx_csr;
  output           pb_cpu_to_io_m1_read_data_valid_sgdma_rx_csr;
  output           pb_cpu_to_io_m1_requests_sgdma_rx_csr;
  output  [  3: 0] sgdma_rx_csr_address;
  output           sgdma_rx_csr_chipselect;
  output           sgdma_rx_csr_irq_from_sa;
  output           sgdma_rx_csr_read;
  output  [ 31: 0] sgdma_rx_csr_readdata_from_sa;
  output           sgdma_rx_csr_reset_n;
  output           sgdma_rx_csr_write;
  output  [ 31: 0] sgdma_rx_csr_writedata;
  input            clk;
  input   [ 22: 0] pb_cpu_to_io_m1_address_to_slave;
  input            pb_cpu_to_io_m1_burstcount;
  input            pb_cpu_to_io_m1_chipselect;
  input            pb_cpu_to_io_m1_latency_counter;
  input            pb_cpu_to_io_m1_read;
  input            pb_cpu_to_io_m1_write;
  input   [ 31: 0] pb_cpu_to_io_m1_writedata;
  input            reset_n;
  input            sgdma_rx_csr_irq;
  input   [ 31: 0] sgdma_rx_csr_readdata;

  reg              d1_reasons_to_wait;
  reg              d1_sgdma_rx_csr_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sgdma_rx_csr;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             pb_cpu_to_io_m1_arbiterlock;
  wire             pb_cpu_to_io_m1_arbiterlock2;
  wire             pb_cpu_to_io_m1_continuerequest;
  wire             pb_cpu_to_io_m1_granted_sgdma_rx_csr;
  wire             pb_cpu_to_io_m1_qualified_request_sgdma_rx_csr;
  wire             pb_cpu_to_io_m1_read_data_valid_sgdma_rx_csr;
  wire             pb_cpu_to_io_m1_requests_sgdma_rx_csr;
  wire             pb_cpu_to_io_m1_saved_grant_sgdma_rx_csr;
  wire    [  3: 0] sgdma_rx_csr_address;
  wire             sgdma_rx_csr_allgrants;
  wire             sgdma_rx_csr_allow_new_arb_cycle;
  wire             sgdma_rx_csr_any_bursting_master_saved_grant;
  wire             sgdma_rx_csr_any_continuerequest;
  wire             sgdma_rx_csr_arb_counter_enable;
  reg              sgdma_rx_csr_arb_share_counter;
  wire             sgdma_rx_csr_arb_share_counter_next_value;
  wire             sgdma_rx_csr_arb_share_set_values;
  wire             sgdma_rx_csr_beginbursttransfer_internal;
  wire             sgdma_rx_csr_begins_xfer;
  wire             sgdma_rx_csr_chipselect;
  wire             sgdma_rx_csr_end_xfer;
  wire             sgdma_rx_csr_firsttransfer;
  wire             sgdma_rx_csr_grant_vector;
  wire             sgdma_rx_csr_in_a_read_cycle;
  wire             sgdma_rx_csr_in_a_write_cycle;
  wire             sgdma_rx_csr_irq_from_sa;
  wire             sgdma_rx_csr_master_qreq_vector;
  wire             sgdma_rx_csr_non_bursting_master_requests;
  wire             sgdma_rx_csr_read;
  wire    [ 31: 0] sgdma_rx_csr_readdata_from_sa;
  reg              sgdma_rx_csr_reg_firsttransfer;
  wire             sgdma_rx_csr_reset_n;
  reg              sgdma_rx_csr_slavearbiterlockenable;
  wire             sgdma_rx_csr_slavearbiterlockenable2;
  wire             sgdma_rx_csr_unreg_firsttransfer;
  wire             sgdma_rx_csr_waits_for_read;
  wire             sgdma_rx_csr_waits_for_write;
  wire             sgdma_rx_csr_write;
  wire    [ 31: 0] sgdma_rx_csr_writedata;
  wire    [ 22: 0] shifted_address_to_sgdma_rx_csr_from_pb_cpu_to_io_m1;
  wire             wait_for_sgdma_rx_csr_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sgdma_rx_csr_end_xfer;
    end


  assign sgdma_rx_csr_begins_xfer = ~d1_reasons_to_wait & ((pb_cpu_to_io_m1_qualified_request_sgdma_rx_csr));
  //assign sgdma_rx_csr_readdata_from_sa = sgdma_rx_csr_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sgdma_rx_csr_readdata_from_sa = sgdma_rx_csr_readdata;

  assign pb_cpu_to_io_m1_requests_sgdma_rx_csr = ({pb_cpu_to_io_m1_address_to_slave[22 : 6] , 6'b0} == 23'h4400) & pb_cpu_to_io_m1_chipselect;
  //sgdma_rx_csr_arb_share_counter set values, which is an e_mux
  assign sgdma_rx_csr_arb_share_set_values = 1;

  //sgdma_rx_csr_non_bursting_master_requests mux, which is an e_mux
  assign sgdma_rx_csr_non_bursting_master_requests = pb_cpu_to_io_m1_requests_sgdma_rx_csr;

  //sgdma_rx_csr_any_bursting_master_saved_grant mux, which is an e_mux
  assign sgdma_rx_csr_any_bursting_master_saved_grant = 0;

  //sgdma_rx_csr_arb_share_counter_next_value assignment, which is an e_assign
  assign sgdma_rx_csr_arb_share_counter_next_value = sgdma_rx_csr_firsttransfer ? (sgdma_rx_csr_arb_share_set_values - 1) : |sgdma_rx_csr_arb_share_counter ? (sgdma_rx_csr_arb_share_counter - 1) : 0;

  //sgdma_rx_csr_allgrants all slave grants, which is an e_mux
  assign sgdma_rx_csr_allgrants = |sgdma_rx_csr_grant_vector;

  //sgdma_rx_csr_end_xfer assignment, which is an e_assign
  assign sgdma_rx_csr_end_xfer = ~(sgdma_rx_csr_waits_for_read | sgdma_rx_csr_waits_for_write);

  //end_xfer_arb_share_counter_term_sgdma_rx_csr arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sgdma_rx_csr = sgdma_rx_csr_end_xfer & (~sgdma_rx_csr_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sgdma_rx_csr_arb_share_counter arbitration counter enable, which is an e_assign
  assign sgdma_rx_csr_arb_counter_enable = (end_xfer_arb_share_counter_term_sgdma_rx_csr & sgdma_rx_csr_allgrants) | (end_xfer_arb_share_counter_term_sgdma_rx_csr & ~sgdma_rx_csr_non_bursting_master_requests);

  //sgdma_rx_csr_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_csr_arb_share_counter <= 0;
      else if (sgdma_rx_csr_arb_counter_enable)
          sgdma_rx_csr_arb_share_counter <= sgdma_rx_csr_arb_share_counter_next_value;
    end


  //sgdma_rx_csr_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_csr_slavearbiterlockenable <= 0;
      else if ((|sgdma_rx_csr_master_qreq_vector & end_xfer_arb_share_counter_term_sgdma_rx_csr) | (end_xfer_arb_share_counter_term_sgdma_rx_csr & ~sgdma_rx_csr_non_bursting_master_requests))
          sgdma_rx_csr_slavearbiterlockenable <= |sgdma_rx_csr_arb_share_counter_next_value;
    end


  //pb_cpu_to_io/m1 sgdma_rx/csr arbiterlock, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock = sgdma_rx_csr_slavearbiterlockenable & pb_cpu_to_io_m1_continuerequest;

  //sgdma_rx_csr_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sgdma_rx_csr_slavearbiterlockenable2 = |sgdma_rx_csr_arb_share_counter_next_value;

  //pb_cpu_to_io/m1 sgdma_rx/csr arbiterlock2, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock2 = sgdma_rx_csr_slavearbiterlockenable2 & pb_cpu_to_io_m1_continuerequest;

  //sgdma_rx_csr_any_continuerequest at least one master continues requesting, which is an e_assign
  assign sgdma_rx_csr_any_continuerequest = 1;

  //pb_cpu_to_io_m1_continuerequest continued request, which is an e_assign
  assign pb_cpu_to_io_m1_continuerequest = 1;

  assign pb_cpu_to_io_m1_qualified_request_sgdma_rx_csr = pb_cpu_to_io_m1_requests_sgdma_rx_csr & ~(((pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ((pb_cpu_to_io_m1_latency_counter != 0))));
  //local readdatavalid pb_cpu_to_io_m1_read_data_valid_sgdma_rx_csr, which is an e_mux
  assign pb_cpu_to_io_m1_read_data_valid_sgdma_rx_csr = pb_cpu_to_io_m1_granted_sgdma_rx_csr & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ~sgdma_rx_csr_waits_for_read;

  //sgdma_rx_csr_writedata mux, which is an e_mux
  assign sgdma_rx_csr_writedata = pb_cpu_to_io_m1_writedata;

  //master is always granted when requested
  assign pb_cpu_to_io_m1_granted_sgdma_rx_csr = pb_cpu_to_io_m1_qualified_request_sgdma_rx_csr;

  //pb_cpu_to_io/m1 saved-grant sgdma_rx/csr, which is an e_assign
  assign pb_cpu_to_io_m1_saved_grant_sgdma_rx_csr = pb_cpu_to_io_m1_requests_sgdma_rx_csr;

  //allow new arb cycle for sgdma_rx/csr, which is an e_assign
  assign sgdma_rx_csr_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign sgdma_rx_csr_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign sgdma_rx_csr_master_qreq_vector = 1;

  //sgdma_rx_csr_reset_n assignment, which is an e_assign
  assign sgdma_rx_csr_reset_n = reset_n;

  assign sgdma_rx_csr_chipselect = pb_cpu_to_io_m1_granted_sgdma_rx_csr;
  //sgdma_rx_csr_firsttransfer first transaction, which is an e_assign
  assign sgdma_rx_csr_firsttransfer = sgdma_rx_csr_begins_xfer ? sgdma_rx_csr_unreg_firsttransfer : sgdma_rx_csr_reg_firsttransfer;

  //sgdma_rx_csr_unreg_firsttransfer first transaction, which is an e_assign
  assign sgdma_rx_csr_unreg_firsttransfer = ~(sgdma_rx_csr_slavearbiterlockenable & sgdma_rx_csr_any_continuerequest);

  //sgdma_rx_csr_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_csr_reg_firsttransfer <= 1'b1;
      else if (sgdma_rx_csr_begins_xfer)
          sgdma_rx_csr_reg_firsttransfer <= sgdma_rx_csr_unreg_firsttransfer;
    end


  //sgdma_rx_csr_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sgdma_rx_csr_beginbursttransfer_internal = sgdma_rx_csr_begins_xfer;

  //sgdma_rx_csr_read assignment, which is an e_mux
  assign sgdma_rx_csr_read = pb_cpu_to_io_m1_granted_sgdma_rx_csr & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect);

  //sgdma_rx_csr_write assignment, which is an e_mux
  assign sgdma_rx_csr_write = pb_cpu_to_io_m1_granted_sgdma_rx_csr & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect);

  assign shifted_address_to_sgdma_rx_csr_from_pb_cpu_to_io_m1 = pb_cpu_to_io_m1_address_to_slave;
  //sgdma_rx_csr_address mux, which is an e_mux
  assign sgdma_rx_csr_address = shifted_address_to_sgdma_rx_csr_from_pb_cpu_to_io_m1 >> 2;

  //d1_sgdma_rx_csr_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sgdma_rx_csr_end_xfer <= 1;
      else 
        d1_sgdma_rx_csr_end_xfer <= sgdma_rx_csr_end_xfer;
    end


  //sgdma_rx_csr_waits_for_read in a cycle, which is an e_mux
  assign sgdma_rx_csr_waits_for_read = sgdma_rx_csr_in_a_read_cycle & sgdma_rx_csr_begins_xfer;

  //sgdma_rx_csr_in_a_read_cycle assignment, which is an e_assign
  assign sgdma_rx_csr_in_a_read_cycle = pb_cpu_to_io_m1_granted_sgdma_rx_csr & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sgdma_rx_csr_in_a_read_cycle;

  //sgdma_rx_csr_waits_for_write in a cycle, which is an e_mux
  assign sgdma_rx_csr_waits_for_write = sgdma_rx_csr_in_a_write_cycle & 0;

  //sgdma_rx_csr_in_a_write_cycle assignment, which is an e_assign
  assign sgdma_rx_csr_in_a_write_cycle = pb_cpu_to_io_m1_granted_sgdma_rx_csr & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sgdma_rx_csr_in_a_write_cycle;

  assign wait_for_sgdma_rx_csr_counter = 0;
  //assign sgdma_rx_csr_irq_from_sa = sgdma_rx_csr_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sgdma_rx_csr_irq_from_sa = sgdma_rx_csr_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_rx/csr enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pb_cpu_to_io/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_io_m1_requests_sgdma_rx_csr && (pb_cpu_to_io_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pb_cpu_to_io/m1 drove 0 on its 'burstcount' port while accessing slave sgdma_rx/csr", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_rx_in_arbitrator (
                                // inputs:
                                 clk,
                                 reset_n,
                                 sgdma_rx_in_ready,
                                 tse_mac_receive_data,
                                 tse_mac_receive_empty,
                                 tse_mac_receive_endofpacket,
                                 tse_mac_receive_error,
                                 tse_mac_receive_startofpacket,
                                 tse_mac_receive_valid,

                                // outputs:
                                 sgdma_rx_in_data,
                                 sgdma_rx_in_empty,
                                 sgdma_rx_in_endofpacket,
                                 sgdma_rx_in_error,
                                 sgdma_rx_in_ready_from_sa,
                                 sgdma_rx_in_startofpacket,
                                 sgdma_rx_in_valid
                              )
;

  output  [ 31: 0] sgdma_rx_in_data;
  output  [  1: 0] sgdma_rx_in_empty;
  output           sgdma_rx_in_endofpacket;
  output  [  5: 0] sgdma_rx_in_error;
  output           sgdma_rx_in_ready_from_sa;
  output           sgdma_rx_in_startofpacket;
  output           sgdma_rx_in_valid;
  input            clk;
  input            reset_n;
  input            sgdma_rx_in_ready;
  input   [ 31: 0] tse_mac_receive_data;
  input   [  1: 0] tse_mac_receive_empty;
  input            tse_mac_receive_endofpacket;
  input   [  5: 0] tse_mac_receive_error;
  input            tse_mac_receive_startofpacket;
  input            tse_mac_receive_valid;

  wire    [ 31: 0] sgdma_rx_in_data;
  wire    [  1: 0] sgdma_rx_in_empty;
  wire             sgdma_rx_in_endofpacket;
  wire    [  5: 0] sgdma_rx_in_error;
  wire             sgdma_rx_in_ready_from_sa;
  wire             sgdma_rx_in_startofpacket;
  wire             sgdma_rx_in_valid;
  //mux sgdma_rx_in_data, which is an e_mux
  assign sgdma_rx_in_data = tse_mac_receive_data;

  //mux sgdma_rx_in_empty, which is an e_mux
  assign sgdma_rx_in_empty = tse_mac_receive_empty;

  //mux sgdma_rx_in_endofpacket, which is an e_mux
  assign sgdma_rx_in_endofpacket = tse_mac_receive_endofpacket;

  //mux sgdma_rx_in_error, which is an e_mux
  assign sgdma_rx_in_error = tse_mac_receive_error;

  //assign sgdma_rx_in_ready_from_sa = sgdma_rx_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sgdma_rx_in_ready_from_sa = sgdma_rx_in_ready;

  //mux sgdma_rx_in_startofpacket, which is an e_mux
  assign sgdma_rx_in_startofpacket = tse_mac_receive_startofpacket;

  //mux sgdma_rx_in_valid, which is an e_mux
  assign sgdma_rx_in_valid = tse_mac_receive_valid;


endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_rx_descriptor_read_arbitrator (
                                             // inputs:
                                              clk,
                                              d1_pb_dma_to_descriptor_memory_s1_end_xfer,
                                              pb_dma_to_descriptor_memory_s1_readdata_from_sa,
                                              pb_dma_to_descriptor_memory_s1_waitrequest_from_sa,
                                              reset_n,
                                              sgdma_rx_descriptor_read_address,
                                              sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1,
                                              sgdma_rx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1,
                                              sgdma_rx_descriptor_read_read,
                                              sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1,
                                              sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register,
                                              sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1,

                                             // outputs:
                                              sgdma_rx_descriptor_read_address_to_slave,
                                              sgdma_rx_descriptor_read_latency_counter,
                                              sgdma_rx_descriptor_read_readdata,
                                              sgdma_rx_descriptor_read_readdatavalid,
                                              sgdma_rx_descriptor_read_waitrequest
                                           )
;

  output  [ 31: 0] sgdma_rx_descriptor_read_address_to_slave;
  output           sgdma_rx_descriptor_read_latency_counter;
  output  [ 31: 0] sgdma_rx_descriptor_read_readdata;
  output           sgdma_rx_descriptor_read_readdatavalid;
  output           sgdma_rx_descriptor_read_waitrequest;
  input            clk;
  input            d1_pb_dma_to_descriptor_memory_s1_end_xfer;
  input   [ 31: 0] pb_dma_to_descriptor_memory_s1_readdata_from_sa;
  input            pb_dma_to_descriptor_memory_s1_waitrequest_from_sa;
  input            reset_n;
  input   [ 31: 0] sgdma_rx_descriptor_read_address;
  input            sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1;
  input            sgdma_rx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1;
  input            sgdma_rx_descriptor_read_read;
  input            sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1;
  input            sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register;
  input            sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_sgdma_rx_descriptor_read_latency_counter;
  wire             pre_flush_sgdma_rx_descriptor_read_readdatavalid;
  wire             r_1;
  reg     [ 31: 0] sgdma_rx_descriptor_read_address_last_time;
  wire    [ 31: 0] sgdma_rx_descriptor_read_address_to_slave;
  wire             sgdma_rx_descriptor_read_is_granted_some_slave;
  reg              sgdma_rx_descriptor_read_latency_counter;
  reg              sgdma_rx_descriptor_read_read_but_no_slave_selected;
  reg              sgdma_rx_descriptor_read_read_last_time;
  wire    [ 31: 0] sgdma_rx_descriptor_read_readdata;
  wire             sgdma_rx_descriptor_read_readdatavalid;
  wire             sgdma_rx_descriptor_read_run;
  wire             sgdma_rx_descriptor_read_waitrequest;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (sgdma_rx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1 | ~sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1) & (sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1 | ~sgdma_rx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1) & ((~sgdma_rx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1 | ~(sgdma_rx_descriptor_read_read) | (1 & ~pb_dma_to_descriptor_memory_s1_waitrequest_from_sa & (sgdma_rx_descriptor_read_read))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_rx_descriptor_read_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_rx_descriptor_read_address_to_slave = {18'b10000000000000,
    sgdma_rx_descriptor_read_address[13 : 0]};

  //sgdma_rx_descriptor_read_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_read_read_but_no_slave_selected <= 0;
      else 
        sgdma_rx_descriptor_read_read_but_no_slave_selected <= sgdma_rx_descriptor_read_read & sgdma_rx_descriptor_read_run & ~sgdma_rx_descriptor_read_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign sgdma_rx_descriptor_read_is_granted_some_slave = sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_sgdma_rx_descriptor_read_readdatavalid = sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign sgdma_rx_descriptor_read_readdatavalid = sgdma_rx_descriptor_read_read_but_no_slave_selected |
    pre_flush_sgdma_rx_descriptor_read_readdatavalid;

  //sgdma_rx/descriptor_read readdata mux, which is an e_mux
  assign sgdma_rx_descriptor_read_readdata = pb_dma_to_descriptor_memory_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign sgdma_rx_descriptor_read_waitrequest = ~sgdma_rx_descriptor_read_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_read_latency_counter <= 0;
      else 
        sgdma_rx_descriptor_read_latency_counter <= p1_sgdma_rx_descriptor_read_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_sgdma_rx_descriptor_read_latency_counter = ((sgdma_rx_descriptor_read_run & sgdma_rx_descriptor_read_read))? latency_load_value :
    (sgdma_rx_descriptor_read_latency_counter)? sgdma_rx_descriptor_read_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_rx_descriptor_read_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_read_address_last_time <= 0;
      else 
        sgdma_rx_descriptor_read_address_last_time <= sgdma_rx_descriptor_read_address;
    end


  //sgdma_rx/descriptor_read waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_rx_descriptor_read_waitrequest & (sgdma_rx_descriptor_read_read);
    end


  //sgdma_rx_descriptor_read_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_descriptor_read_address != sgdma_rx_descriptor_read_address_last_time))
        begin
          $write("%0d ns: sgdma_rx_descriptor_read_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_descriptor_read_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_read_read_last_time <= 0;
      else 
        sgdma_rx_descriptor_read_read_last_time <= sgdma_rx_descriptor_read_read;
    end


  //sgdma_rx_descriptor_read_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_descriptor_read_read != sgdma_rx_descriptor_read_read_last_time))
        begin
          $write("%0d ns: sgdma_rx_descriptor_read_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_rx_descriptor_write_arbitrator (
                                              // inputs:
                                               clk,
                                               d1_pb_dma_to_descriptor_memory_s1_end_xfer,
                                               pb_dma_to_descriptor_memory_s1_waitrequest_from_sa,
                                               reset_n,
                                               sgdma_rx_descriptor_write_address,
                                               sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1,
                                               sgdma_rx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1,
                                               sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1,
                                               sgdma_rx_descriptor_write_write,
                                               sgdma_rx_descriptor_write_writedata,

                                              // outputs:
                                               sgdma_rx_descriptor_write_address_to_slave,
                                               sgdma_rx_descriptor_write_waitrequest
                                            )
;

  output  [ 31: 0] sgdma_rx_descriptor_write_address_to_slave;
  output           sgdma_rx_descriptor_write_waitrequest;
  input            clk;
  input            d1_pb_dma_to_descriptor_memory_s1_end_xfer;
  input            pb_dma_to_descriptor_memory_s1_waitrequest_from_sa;
  input            reset_n;
  input   [ 31: 0] sgdma_rx_descriptor_write_address;
  input            sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1;
  input            sgdma_rx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1;
  input            sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1;
  input            sgdma_rx_descriptor_write_write;
  input   [ 31: 0] sgdma_rx_descriptor_write_writedata;

  reg              active_and_waiting_last_time;
  wire             r_1;
  reg     [ 31: 0] sgdma_rx_descriptor_write_address_last_time;
  wire    [ 31: 0] sgdma_rx_descriptor_write_address_to_slave;
  wire             sgdma_rx_descriptor_write_run;
  wire             sgdma_rx_descriptor_write_waitrequest;
  reg              sgdma_rx_descriptor_write_write_last_time;
  reg     [ 31: 0] sgdma_rx_descriptor_write_writedata_last_time;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (sgdma_rx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1 | ~sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1) & (sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1 | ~sgdma_rx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1) & ((~sgdma_rx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1 | ~(sgdma_rx_descriptor_write_write) | (1 & ~pb_dma_to_descriptor_memory_s1_waitrequest_from_sa & (sgdma_rx_descriptor_write_write))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_rx_descriptor_write_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_rx_descriptor_write_address_to_slave = {18'b10000000000000,
    sgdma_rx_descriptor_write_address[13 : 0]};

  //actual waitrequest port, which is an e_assign
  assign sgdma_rx_descriptor_write_waitrequest = ~sgdma_rx_descriptor_write_run;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_rx_descriptor_write_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_write_address_last_time <= 0;
      else 
        sgdma_rx_descriptor_write_address_last_time <= sgdma_rx_descriptor_write_address;
    end


  //sgdma_rx/descriptor_write waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_rx_descriptor_write_waitrequest & (sgdma_rx_descriptor_write_write);
    end


  //sgdma_rx_descriptor_write_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_descriptor_write_address != sgdma_rx_descriptor_write_address_last_time))
        begin
          $write("%0d ns: sgdma_rx_descriptor_write_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_descriptor_write_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_write_write_last_time <= 0;
      else 
        sgdma_rx_descriptor_write_write_last_time <= sgdma_rx_descriptor_write_write;
    end


  //sgdma_rx_descriptor_write_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_descriptor_write_write != sgdma_rx_descriptor_write_write_last_time))
        begin
          $write("%0d ns: sgdma_rx_descriptor_write_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_descriptor_write_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_write_writedata_last_time <= 0;
      else 
        sgdma_rx_descriptor_write_writedata_last_time <= sgdma_rx_descriptor_write_writedata;
    end


  //sgdma_rx_descriptor_write_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_descriptor_write_writedata != sgdma_rx_descriptor_write_writedata_last_time) & sgdma_rx_descriptor_write_write)
        begin
          $write("%0d ns: sgdma_rx_descriptor_write_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_rx_m_write_arbitrator (
                                     // inputs:
                                      clk,
                                      d1_pb_dma_to_ddr3_top_s1_end_xfer,
                                      pb_dma_to_ddr3_top_s1_waitrequest_from_sa,
                                      reset_n,
                                      sgdma_rx_m_write_address,
                                      sgdma_rx_m_write_byteenable,
                                      sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1,
                                      sgdma_rx_m_write_qualified_request_pb_dma_to_ddr3_top_s1,
                                      sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1,
                                      sgdma_rx_m_write_write,
                                      sgdma_rx_m_write_writedata,

                                     // outputs:
                                      sgdma_rx_m_write_address_to_slave,
                                      sgdma_rx_m_write_waitrequest
                                   )
;

  output  [ 31: 0] sgdma_rx_m_write_address_to_slave;
  output           sgdma_rx_m_write_waitrequest;
  input            clk;
  input            d1_pb_dma_to_ddr3_top_s1_end_xfer;
  input            pb_dma_to_ddr3_top_s1_waitrequest_from_sa;
  input            reset_n;
  input   [ 31: 0] sgdma_rx_m_write_address;
  input   [  3: 0] sgdma_rx_m_write_byteenable;
  input            sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1;
  input            sgdma_rx_m_write_qualified_request_pb_dma_to_ddr3_top_s1;
  input            sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1;
  input            sgdma_rx_m_write_write;
  input   [ 31: 0] sgdma_rx_m_write_writedata;

  reg              active_and_waiting_last_time;
  wire             r_1;
  reg     [ 31: 0] sgdma_rx_m_write_address_last_time;
  wire    [ 31: 0] sgdma_rx_m_write_address_to_slave;
  reg     [  3: 0] sgdma_rx_m_write_byteenable_last_time;
  wire             sgdma_rx_m_write_run;
  wire             sgdma_rx_m_write_waitrequest;
  reg              sgdma_rx_m_write_write_last_time;
  reg     [ 31: 0] sgdma_rx_m_write_writedata_last_time;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (sgdma_rx_m_write_qualified_request_pb_dma_to_ddr3_top_s1 | ~sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1) & (sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1 | ~sgdma_rx_m_write_qualified_request_pb_dma_to_ddr3_top_s1) & ((~sgdma_rx_m_write_qualified_request_pb_dma_to_ddr3_top_s1 | ~(sgdma_rx_m_write_write) | (1 & ~pb_dma_to_ddr3_top_s1_waitrequest_from_sa & (sgdma_rx_m_write_write))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_rx_m_write_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_rx_m_write_address_to_slave = {5'b10,
    sgdma_rx_m_write_address[26 : 0]};

  //actual waitrequest port, which is an e_assign
  assign sgdma_rx_m_write_waitrequest = ~sgdma_rx_m_write_run;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_rx_m_write_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_m_write_address_last_time <= 0;
      else 
        sgdma_rx_m_write_address_last_time <= sgdma_rx_m_write_address;
    end


  //sgdma_rx/m_write waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_rx_m_write_waitrequest & (sgdma_rx_m_write_write);
    end


  //sgdma_rx_m_write_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_m_write_address != sgdma_rx_m_write_address_last_time))
        begin
          $write("%0d ns: sgdma_rx_m_write_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_m_write_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_m_write_byteenable_last_time <= 0;
      else 
        sgdma_rx_m_write_byteenable_last_time <= sgdma_rx_m_write_byteenable;
    end


  //sgdma_rx_m_write_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_m_write_byteenable != sgdma_rx_m_write_byteenable_last_time))
        begin
          $write("%0d ns: sgdma_rx_m_write_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_m_write_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_m_write_write_last_time <= 0;
      else 
        sgdma_rx_m_write_write_last_time <= sgdma_rx_m_write_write;
    end


  //sgdma_rx_m_write_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_m_write_write != sgdma_rx_m_write_write_last_time))
        begin
          $write("%0d ns: sgdma_rx_m_write_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_m_write_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_m_write_writedata_last_time <= 0;
      else 
        sgdma_rx_m_write_writedata_last_time <= sgdma_rx_m_write_writedata;
    end


  //sgdma_rx_m_write_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_m_write_writedata != sgdma_rx_m_write_writedata_last_time) & sgdma_rx_m_write_write)
        begin
          $write("%0d ns: sgdma_rx_m_write_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_tx_csr_arbitrator (
                                 // inputs:
                                  clk,
                                  pb_cpu_to_io_m1_address_to_slave,
                                  pb_cpu_to_io_m1_burstcount,
                                  pb_cpu_to_io_m1_chipselect,
                                  pb_cpu_to_io_m1_latency_counter,
                                  pb_cpu_to_io_m1_read,
                                  pb_cpu_to_io_m1_write,
                                  pb_cpu_to_io_m1_writedata,
                                  reset_n,
                                  sgdma_tx_csr_irq,
                                  sgdma_tx_csr_readdata,

                                 // outputs:
                                  d1_sgdma_tx_csr_end_xfer,
                                  pb_cpu_to_io_m1_granted_sgdma_tx_csr,
                                  pb_cpu_to_io_m1_qualified_request_sgdma_tx_csr,
                                  pb_cpu_to_io_m1_read_data_valid_sgdma_tx_csr,
                                  pb_cpu_to_io_m1_requests_sgdma_tx_csr,
                                  sgdma_tx_csr_address,
                                  sgdma_tx_csr_chipselect,
                                  sgdma_tx_csr_irq_from_sa,
                                  sgdma_tx_csr_read,
                                  sgdma_tx_csr_readdata_from_sa,
                                  sgdma_tx_csr_reset_n,
                                  sgdma_tx_csr_write,
                                  sgdma_tx_csr_writedata
                               )
;

  output           d1_sgdma_tx_csr_end_xfer;
  output           pb_cpu_to_io_m1_granted_sgdma_tx_csr;
  output           pb_cpu_to_io_m1_qualified_request_sgdma_tx_csr;
  output           pb_cpu_to_io_m1_read_data_valid_sgdma_tx_csr;
  output           pb_cpu_to_io_m1_requests_sgdma_tx_csr;
  output  [  3: 0] sgdma_tx_csr_address;
  output           sgdma_tx_csr_chipselect;
  output           sgdma_tx_csr_irq_from_sa;
  output           sgdma_tx_csr_read;
  output  [ 31: 0] sgdma_tx_csr_readdata_from_sa;
  output           sgdma_tx_csr_reset_n;
  output           sgdma_tx_csr_write;
  output  [ 31: 0] sgdma_tx_csr_writedata;
  input            clk;
  input   [ 22: 0] pb_cpu_to_io_m1_address_to_slave;
  input            pb_cpu_to_io_m1_burstcount;
  input            pb_cpu_to_io_m1_chipselect;
  input            pb_cpu_to_io_m1_latency_counter;
  input            pb_cpu_to_io_m1_read;
  input            pb_cpu_to_io_m1_write;
  input   [ 31: 0] pb_cpu_to_io_m1_writedata;
  input            reset_n;
  input            sgdma_tx_csr_irq;
  input   [ 31: 0] sgdma_tx_csr_readdata;

  reg              d1_reasons_to_wait;
  reg              d1_sgdma_tx_csr_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sgdma_tx_csr;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             pb_cpu_to_io_m1_arbiterlock;
  wire             pb_cpu_to_io_m1_arbiterlock2;
  wire             pb_cpu_to_io_m1_continuerequest;
  wire             pb_cpu_to_io_m1_granted_sgdma_tx_csr;
  wire             pb_cpu_to_io_m1_qualified_request_sgdma_tx_csr;
  wire             pb_cpu_to_io_m1_read_data_valid_sgdma_tx_csr;
  wire             pb_cpu_to_io_m1_requests_sgdma_tx_csr;
  wire             pb_cpu_to_io_m1_saved_grant_sgdma_tx_csr;
  wire    [  3: 0] sgdma_tx_csr_address;
  wire             sgdma_tx_csr_allgrants;
  wire             sgdma_tx_csr_allow_new_arb_cycle;
  wire             sgdma_tx_csr_any_bursting_master_saved_grant;
  wire             sgdma_tx_csr_any_continuerequest;
  wire             sgdma_tx_csr_arb_counter_enable;
  reg              sgdma_tx_csr_arb_share_counter;
  wire             sgdma_tx_csr_arb_share_counter_next_value;
  wire             sgdma_tx_csr_arb_share_set_values;
  wire             sgdma_tx_csr_beginbursttransfer_internal;
  wire             sgdma_tx_csr_begins_xfer;
  wire             sgdma_tx_csr_chipselect;
  wire             sgdma_tx_csr_end_xfer;
  wire             sgdma_tx_csr_firsttransfer;
  wire             sgdma_tx_csr_grant_vector;
  wire             sgdma_tx_csr_in_a_read_cycle;
  wire             sgdma_tx_csr_in_a_write_cycle;
  wire             sgdma_tx_csr_irq_from_sa;
  wire             sgdma_tx_csr_master_qreq_vector;
  wire             sgdma_tx_csr_non_bursting_master_requests;
  wire             sgdma_tx_csr_read;
  wire    [ 31: 0] sgdma_tx_csr_readdata_from_sa;
  reg              sgdma_tx_csr_reg_firsttransfer;
  wire             sgdma_tx_csr_reset_n;
  reg              sgdma_tx_csr_slavearbiterlockenable;
  wire             sgdma_tx_csr_slavearbiterlockenable2;
  wire             sgdma_tx_csr_unreg_firsttransfer;
  wire             sgdma_tx_csr_waits_for_read;
  wire             sgdma_tx_csr_waits_for_write;
  wire             sgdma_tx_csr_write;
  wire    [ 31: 0] sgdma_tx_csr_writedata;
  wire    [ 22: 0] shifted_address_to_sgdma_tx_csr_from_pb_cpu_to_io_m1;
  wire             wait_for_sgdma_tx_csr_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sgdma_tx_csr_end_xfer;
    end


  assign sgdma_tx_csr_begins_xfer = ~d1_reasons_to_wait & ((pb_cpu_to_io_m1_qualified_request_sgdma_tx_csr));
  //assign sgdma_tx_csr_readdata_from_sa = sgdma_tx_csr_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sgdma_tx_csr_readdata_from_sa = sgdma_tx_csr_readdata;

  assign pb_cpu_to_io_m1_requests_sgdma_tx_csr = ({pb_cpu_to_io_m1_address_to_slave[22 : 6] , 6'b0} == 23'h4800) & pb_cpu_to_io_m1_chipselect;
  //sgdma_tx_csr_arb_share_counter set values, which is an e_mux
  assign sgdma_tx_csr_arb_share_set_values = 1;

  //sgdma_tx_csr_non_bursting_master_requests mux, which is an e_mux
  assign sgdma_tx_csr_non_bursting_master_requests = pb_cpu_to_io_m1_requests_sgdma_tx_csr;

  //sgdma_tx_csr_any_bursting_master_saved_grant mux, which is an e_mux
  assign sgdma_tx_csr_any_bursting_master_saved_grant = 0;

  //sgdma_tx_csr_arb_share_counter_next_value assignment, which is an e_assign
  assign sgdma_tx_csr_arb_share_counter_next_value = sgdma_tx_csr_firsttransfer ? (sgdma_tx_csr_arb_share_set_values - 1) : |sgdma_tx_csr_arb_share_counter ? (sgdma_tx_csr_arb_share_counter - 1) : 0;

  //sgdma_tx_csr_allgrants all slave grants, which is an e_mux
  assign sgdma_tx_csr_allgrants = |sgdma_tx_csr_grant_vector;

  //sgdma_tx_csr_end_xfer assignment, which is an e_assign
  assign sgdma_tx_csr_end_xfer = ~(sgdma_tx_csr_waits_for_read | sgdma_tx_csr_waits_for_write);

  //end_xfer_arb_share_counter_term_sgdma_tx_csr arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sgdma_tx_csr = sgdma_tx_csr_end_xfer & (~sgdma_tx_csr_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sgdma_tx_csr_arb_share_counter arbitration counter enable, which is an e_assign
  assign sgdma_tx_csr_arb_counter_enable = (end_xfer_arb_share_counter_term_sgdma_tx_csr & sgdma_tx_csr_allgrants) | (end_xfer_arb_share_counter_term_sgdma_tx_csr & ~sgdma_tx_csr_non_bursting_master_requests);

  //sgdma_tx_csr_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_csr_arb_share_counter <= 0;
      else if (sgdma_tx_csr_arb_counter_enable)
          sgdma_tx_csr_arb_share_counter <= sgdma_tx_csr_arb_share_counter_next_value;
    end


  //sgdma_tx_csr_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_csr_slavearbiterlockenable <= 0;
      else if ((|sgdma_tx_csr_master_qreq_vector & end_xfer_arb_share_counter_term_sgdma_tx_csr) | (end_xfer_arb_share_counter_term_sgdma_tx_csr & ~sgdma_tx_csr_non_bursting_master_requests))
          sgdma_tx_csr_slavearbiterlockenable <= |sgdma_tx_csr_arb_share_counter_next_value;
    end


  //pb_cpu_to_io/m1 sgdma_tx/csr arbiterlock, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock = sgdma_tx_csr_slavearbiterlockenable & pb_cpu_to_io_m1_continuerequest;

  //sgdma_tx_csr_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sgdma_tx_csr_slavearbiterlockenable2 = |sgdma_tx_csr_arb_share_counter_next_value;

  //pb_cpu_to_io/m1 sgdma_tx/csr arbiterlock2, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock2 = sgdma_tx_csr_slavearbiterlockenable2 & pb_cpu_to_io_m1_continuerequest;

  //sgdma_tx_csr_any_continuerequest at least one master continues requesting, which is an e_assign
  assign sgdma_tx_csr_any_continuerequest = 1;

  //pb_cpu_to_io_m1_continuerequest continued request, which is an e_assign
  assign pb_cpu_to_io_m1_continuerequest = 1;

  assign pb_cpu_to_io_m1_qualified_request_sgdma_tx_csr = pb_cpu_to_io_m1_requests_sgdma_tx_csr & ~(((pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ((pb_cpu_to_io_m1_latency_counter != 0))));
  //local readdatavalid pb_cpu_to_io_m1_read_data_valid_sgdma_tx_csr, which is an e_mux
  assign pb_cpu_to_io_m1_read_data_valid_sgdma_tx_csr = pb_cpu_to_io_m1_granted_sgdma_tx_csr & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ~sgdma_tx_csr_waits_for_read;

  //sgdma_tx_csr_writedata mux, which is an e_mux
  assign sgdma_tx_csr_writedata = pb_cpu_to_io_m1_writedata;

  //master is always granted when requested
  assign pb_cpu_to_io_m1_granted_sgdma_tx_csr = pb_cpu_to_io_m1_qualified_request_sgdma_tx_csr;

  //pb_cpu_to_io/m1 saved-grant sgdma_tx/csr, which is an e_assign
  assign pb_cpu_to_io_m1_saved_grant_sgdma_tx_csr = pb_cpu_to_io_m1_requests_sgdma_tx_csr;

  //allow new arb cycle for sgdma_tx/csr, which is an e_assign
  assign sgdma_tx_csr_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign sgdma_tx_csr_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign sgdma_tx_csr_master_qreq_vector = 1;

  //sgdma_tx_csr_reset_n assignment, which is an e_assign
  assign sgdma_tx_csr_reset_n = reset_n;

  assign sgdma_tx_csr_chipselect = pb_cpu_to_io_m1_granted_sgdma_tx_csr;
  //sgdma_tx_csr_firsttransfer first transaction, which is an e_assign
  assign sgdma_tx_csr_firsttransfer = sgdma_tx_csr_begins_xfer ? sgdma_tx_csr_unreg_firsttransfer : sgdma_tx_csr_reg_firsttransfer;

  //sgdma_tx_csr_unreg_firsttransfer first transaction, which is an e_assign
  assign sgdma_tx_csr_unreg_firsttransfer = ~(sgdma_tx_csr_slavearbiterlockenable & sgdma_tx_csr_any_continuerequest);

  //sgdma_tx_csr_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_csr_reg_firsttransfer <= 1'b1;
      else if (sgdma_tx_csr_begins_xfer)
          sgdma_tx_csr_reg_firsttransfer <= sgdma_tx_csr_unreg_firsttransfer;
    end


  //sgdma_tx_csr_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sgdma_tx_csr_beginbursttransfer_internal = sgdma_tx_csr_begins_xfer;

  //sgdma_tx_csr_read assignment, which is an e_mux
  assign sgdma_tx_csr_read = pb_cpu_to_io_m1_granted_sgdma_tx_csr & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect);

  //sgdma_tx_csr_write assignment, which is an e_mux
  assign sgdma_tx_csr_write = pb_cpu_to_io_m1_granted_sgdma_tx_csr & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect);

  assign shifted_address_to_sgdma_tx_csr_from_pb_cpu_to_io_m1 = pb_cpu_to_io_m1_address_to_slave;
  //sgdma_tx_csr_address mux, which is an e_mux
  assign sgdma_tx_csr_address = shifted_address_to_sgdma_tx_csr_from_pb_cpu_to_io_m1 >> 2;

  //d1_sgdma_tx_csr_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sgdma_tx_csr_end_xfer <= 1;
      else 
        d1_sgdma_tx_csr_end_xfer <= sgdma_tx_csr_end_xfer;
    end


  //sgdma_tx_csr_waits_for_read in a cycle, which is an e_mux
  assign sgdma_tx_csr_waits_for_read = sgdma_tx_csr_in_a_read_cycle & sgdma_tx_csr_begins_xfer;

  //sgdma_tx_csr_in_a_read_cycle assignment, which is an e_assign
  assign sgdma_tx_csr_in_a_read_cycle = pb_cpu_to_io_m1_granted_sgdma_tx_csr & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sgdma_tx_csr_in_a_read_cycle;

  //sgdma_tx_csr_waits_for_write in a cycle, which is an e_mux
  assign sgdma_tx_csr_waits_for_write = sgdma_tx_csr_in_a_write_cycle & 0;

  //sgdma_tx_csr_in_a_write_cycle assignment, which is an e_assign
  assign sgdma_tx_csr_in_a_write_cycle = pb_cpu_to_io_m1_granted_sgdma_tx_csr & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sgdma_tx_csr_in_a_write_cycle;

  assign wait_for_sgdma_tx_csr_counter = 0;
  //assign sgdma_tx_csr_irq_from_sa = sgdma_tx_csr_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sgdma_tx_csr_irq_from_sa = sgdma_tx_csr_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_tx/csr enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pb_cpu_to_io/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_io_m1_requests_sgdma_tx_csr && (pb_cpu_to_io_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pb_cpu_to_io/m1 drove 0 on its 'burstcount' port while accessing slave sgdma_tx/csr", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_tx_descriptor_read_arbitrator (
                                             // inputs:
                                              clk,
                                              d1_pb_dma_to_descriptor_memory_s1_end_xfer,
                                              pb_dma_to_descriptor_memory_s1_readdata_from_sa,
                                              pb_dma_to_descriptor_memory_s1_waitrequest_from_sa,
                                              reset_n,
                                              sgdma_tx_descriptor_read_address,
                                              sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1,
                                              sgdma_tx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1,
                                              sgdma_tx_descriptor_read_read,
                                              sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1,
                                              sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register,
                                              sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1,

                                             // outputs:
                                              sgdma_tx_descriptor_read_address_to_slave,
                                              sgdma_tx_descriptor_read_latency_counter,
                                              sgdma_tx_descriptor_read_readdata,
                                              sgdma_tx_descriptor_read_readdatavalid,
                                              sgdma_tx_descriptor_read_waitrequest
                                           )
;

  output  [ 31: 0] sgdma_tx_descriptor_read_address_to_slave;
  output           sgdma_tx_descriptor_read_latency_counter;
  output  [ 31: 0] sgdma_tx_descriptor_read_readdata;
  output           sgdma_tx_descriptor_read_readdatavalid;
  output           sgdma_tx_descriptor_read_waitrequest;
  input            clk;
  input            d1_pb_dma_to_descriptor_memory_s1_end_xfer;
  input   [ 31: 0] pb_dma_to_descriptor_memory_s1_readdata_from_sa;
  input            pb_dma_to_descriptor_memory_s1_waitrequest_from_sa;
  input            reset_n;
  input   [ 31: 0] sgdma_tx_descriptor_read_address;
  input            sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1;
  input            sgdma_tx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1;
  input            sgdma_tx_descriptor_read_read;
  input            sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1;
  input            sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register;
  input            sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_sgdma_tx_descriptor_read_latency_counter;
  wire             pre_flush_sgdma_tx_descriptor_read_readdatavalid;
  wire             r_1;
  reg     [ 31: 0] sgdma_tx_descriptor_read_address_last_time;
  wire    [ 31: 0] sgdma_tx_descriptor_read_address_to_slave;
  wire             sgdma_tx_descriptor_read_is_granted_some_slave;
  reg              sgdma_tx_descriptor_read_latency_counter;
  reg              sgdma_tx_descriptor_read_read_but_no_slave_selected;
  reg              sgdma_tx_descriptor_read_read_last_time;
  wire    [ 31: 0] sgdma_tx_descriptor_read_readdata;
  wire             sgdma_tx_descriptor_read_readdatavalid;
  wire             sgdma_tx_descriptor_read_run;
  wire             sgdma_tx_descriptor_read_waitrequest;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (sgdma_tx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1 | ~sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1) & (sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1 | ~sgdma_tx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1) & ((~sgdma_tx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1 | ~(sgdma_tx_descriptor_read_read) | (1 & ~pb_dma_to_descriptor_memory_s1_waitrequest_from_sa & (sgdma_tx_descriptor_read_read))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_tx_descriptor_read_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_tx_descriptor_read_address_to_slave = {18'b10000000000000,
    sgdma_tx_descriptor_read_address[13 : 0]};

  //sgdma_tx_descriptor_read_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_read_read_but_no_slave_selected <= 0;
      else 
        sgdma_tx_descriptor_read_read_but_no_slave_selected <= sgdma_tx_descriptor_read_read & sgdma_tx_descriptor_read_run & ~sgdma_tx_descriptor_read_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign sgdma_tx_descriptor_read_is_granted_some_slave = sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_sgdma_tx_descriptor_read_readdatavalid = sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign sgdma_tx_descriptor_read_readdatavalid = sgdma_tx_descriptor_read_read_but_no_slave_selected |
    pre_flush_sgdma_tx_descriptor_read_readdatavalid;

  //sgdma_tx/descriptor_read readdata mux, which is an e_mux
  assign sgdma_tx_descriptor_read_readdata = pb_dma_to_descriptor_memory_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign sgdma_tx_descriptor_read_waitrequest = ~sgdma_tx_descriptor_read_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_read_latency_counter <= 0;
      else 
        sgdma_tx_descriptor_read_latency_counter <= p1_sgdma_tx_descriptor_read_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_sgdma_tx_descriptor_read_latency_counter = ((sgdma_tx_descriptor_read_run & sgdma_tx_descriptor_read_read))? latency_load_value :
    (sgdma_tx_descriptor_read_latency_counter)? sgdma_tx_descriptor_read_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_tx_descriptor_read_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_read_address_last_time <= 0;
      else 
        sgdma_tx_descriptor_read_address_last_time <= sgdma_tx_descriptor_read_address;
    end


  //sgdma_tx/descriptor_read waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_tx_descriptor_read_waitrequest & (sgdma_tx_descriptor_read_read);
    end


  //sgdma_tx_descriptor_read_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_descriptor_read_address != sgdma_tx_descriptor_read_address_last_time))
        begin
          $write("%0d ns: sgdma_tx_descriptor_read_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_tx_descriptor_read_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_read_read_last_time <= 0;
      else 
        sgdma_tx_descriptor_read_read_last_time <= sgdma_tx_descriptor_read_read;
    end


  //sgdma_tx_descriptor_read_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_descriptor_read_read != sgdma_tx_descriptor_read_read_last_time))
        begin
          $write("%0d ns: sgdma_tx_descriptor_read_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_tx_descriptor_write_arbitrator (
                                              // inputs:
                                               clk,
                                               d1_pb_dma_to_descriptor_memory_s1_end_xfer,
                                               pb_dma_to_descriptor_memory_s1_waitrequest_from_sa,
                                               reset_n,
                                               sgdma_tx_descriptor_write_address,
                                               sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1,
                                               sgdma_tx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1,
                                               sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1,
                                               sgdma_tx_descriptor_write_write,
                                               sgdma_tx_descriptor_write_writedata,

                                              // outputs:
                                               sgdma_tx_descriptor_write_address_to_slave,
                                               sgdma_tx_descriptor_write_waitrequest
                                            )
;

  output  [ 31: 0] sgdma_tx_descriptor_write_address_to_slave;
  output           sgdma_tx_descriptor_write_waitrequest;
  input            clk;
  input            d1_pb_dma_to_descriptor_memory_s1_end_xfer;
  input            pb_dma_to_descriptor_memory_s1_waitrequest_from_sa;
  input            reset_n;
  input   [ 31: 0] sgdma_tx_descriptor_write_address;
  input            sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1;
  input            sgdma_tx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1;
  input            sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1;
  input            sgdma_tx_descriptor_write_write;
  input   [ 31: 0] sgdma_tx_descriptor_write_writedata;

  reg              active_and_waiting_last_time;
  wire             r_1;
  reg     [ 31: 0] sgdma_tx_descriptor_write_address_last_time;
  wire    [ 31: 0] sgdma_tx_descriptor_write_address_to_slave;
  wire             sgdma_tx_descriptor_write_run;
  wire             sgdma_tx_descriptor_write_waitrequest;
  reg              sgdma_tx_descriptor_write_write_last_time;
  reg     [ 31: 0] sgdma_tx_descriptor_write_writedata_last_time;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (sgdma_tx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1 | ~sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1) & (sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1 | ~sgdma_tx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1) & ((~sgdma_tx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1 | ~(sgdma_tx_descriptor_write_write) | (1 & ~pb_dma_to_descriptor_memory_s1_waitrequest_from_sa & (sgdma_tx_descriptor_write_write))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_tx_descriptor_write_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_tx_descriptor_write_address_to_slave = {18'b10000000000000,
    sgdma_tx_descriptor_write_address[13 : 0]};

  //actual waitrequest port, which is an e_assign
  assign sgdma_tx_descriptor_write_waitrequest = ~sgdma_tx_descriptor_write_run;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_tx_descriptor_write_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_write_address_last_time <= 0;
      else 
        sgdma_tx_descriptor_write_address_last_time <= sgdma_tx_descriptor_write_address;
    end


  //sgdma_tx/descriptor_write waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_tx_descriptor_write_waitrequest & (sgdma_tx_descriptor_write_write);
    end


  //sgdma_tx_descriptor_write_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_descriptor_write_address != sgdma_tx_descriptor_write_address_last_time))
        begin
          $write("%0d ns: sgdma_tx_descriptor_write_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_tx_descriptor_write_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_write_write_last_time <= 0;
      else 
        sgdma_tx_descriptor_write_write_last_time <= sgdma_tx_descriptor_write_write;
    end


  //sgdma_tx_descriptor_write_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_descriptor_write_write != sgdma_tx_descriptor_write_write_last_time))
        begin
          $write("%0d ns: sgdma_tx_descriptor_write_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_tx_descriptor_write_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_write_writedata_last_time <= 0;
      else 
        sgdma_tx_descriptor_write_writedata_last_time <= sgdma_tx_descriptor_write_writedata;
    end


  //sgdma_tx_descriptor_write_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_descriptor_write_writedata != sgdma_tx_descriptor_write_writedata_last_time) & sgdma_tx_descriptor_write_write)
        begin
          $write("%0d ns: sgdma_tx_descriptor_write_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_tx_m_read_arbitrator (
                                    // inputs:
                                     clk,
                                     d1_pb_dma_to_ddr3_top_s1_end_xfer,
                                     pb_dma_to_ddr3_top_s1_readdata_from_sa,
                                     pb_dma_to_ddr3_top_s1_waitrequest_from_sa,
                                     reset_n,
                                     sgdma_tx_m_read_address,
                                     sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1,
                                     sgdma_tx_m_read_qualified_request_pb_dma_to_ddr3_top_s1,
                                     sgdma_tx_m_read_read,
                                     sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1,
                                     sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1_shift_register,
                                     sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1,

                                    // outputs:
                                     sgdma_tx_m_read_address_to_slave,
                                     sgdma_tx_m_read_latency_counter,
                                     sgdma_tx_m_read_readdata,
                                     sgdma_tx_m_read_readdatavalid,
                                     sgdma_tx_m_read_waitrequest
                                  )
;

  output  [ 31: 0] sgdma_tx_m_read_address_to_slave;
  output           sgdma_tx_m_read_latency_counter;
  output  [ 31: 0] sgdma_tx_m_read_readdata;
  output           sgdma_tx_m_read_readdatavalid;
  output           sgdma_tx_m_read_waitrequest;
  input            clk;
  input            d1_pb_dma_to_ddr3_top_s1_end_xfer;
  input   [ 31: 0] pb_dma_to_ddr3_top_s1_readdata_from_sa;
  input            pb_dma_to_ddr3_top_s1_waitrequest_from_sa;
  input            reset_n;
  input   [ 31: 0] sgdma_tx_m_read_address;
  input            sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1;
  input            sgdma_tx_m_read_qualified_request_pb_dma_to_ddr3_top_s1;
  input            sgdma_tx_m_read_read;
  input            sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1;
  input            sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1_shift_register;
  input            sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_sgdma_tx_m_read_latency_counter;
  wire             pre_flush_sgdma_tx_m_read_readdatavalid;
  wire             r_1;
  reg     [ 31: 0] sgdma_tx_m_read_address_last_time;
  wire    [ 31: 0] sgdma_tx_m_read_address_to_slave;
  wire             sgdma_tx_m_read_is_granted_some_slave;
  reg              sgdma_tx_m_read_latency_counter;
  reg              sgdma_tx_m_read_read_but_no_slave_selected;
  reg              sgdma_tx_m_read_read_last_time;
  wire    [ 31: 0] sgdma_tx_m_read_readdata;
  wire             sgdma_tx_m_read_readdatavalid;
  wire             sgdma_tx_m_read_run;
  wire             sgdma_tx_m_read_waitrequest;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (sgdma_tx_m_read_qualified_request_pb_dma_to_ddr3_top_s1 | ~sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1) & (sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1 | ~sgdma_tx_m_read_qualified_request_pb_dma_to_ddr3_top_s1) & ((~sgdma_tx_m_read_qualified_request_pb_dma_to_ddr3_top_s1 | ~(sgdma_tx_m_read_read) | (1 & ~pb_dma_to_ddr3_top_s1_waitrequest_from_sa & (sgdma_tx_m_read_read))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_tx_m_read_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_tx_m_read_address_to_slave = {5'b10,
    sgdma_tx_m_read_address[26 : 0]};

  //sgdma_tx_m_read_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_m_read_read_but_no_slave_selected <= 0;
      else 
        sgdma_tx_m_read_read_but_no_slave_selected <= sgdma_tx_m_read_read & sgdma_tx_m_read_run & ~sgdma_tx_m_read_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign sgdma_tx_m_read_is_granted_some_slave = sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_sgdma_tx_m_read_readdatavalid = sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign sgdma_tx_m_read_readdatavalid = sgdma_tx_m_read_read_but_no_slave_selected |
    pre_flush_sgdma_tx_m_read_readdatavalid;

  //sgdma_tx/m_read readdata mux, which is an e_mux
  assign sgdma_tx_m_read_readdata = pb_dma_to_ddr3_top_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign sgdma_tx_m_read_waitrequest = ~sgdma_tx_m_read_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_m_read_latency_counter <= 0;
      else 
        sgdma_tx_m_read_latency_counter <= p1_sgdma_tx_m_read_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_sgdma_tx_m_read_latency_counter = ((sgdma_tx_m_read_run & sgdma_tx_m_read_read))? latency_load_value :
    (sgdma_tx_m_read_latency_counter)? sgdma_tx_m_read_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_tx_m_read_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_m_read_address_last_time <= 0;
      else 
        sgdma_tx_m_read_address_last_time <= sgdma_tx_m_read_address;
    end


  //sgdma_tx/m_read waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_tx_m_read_waitrequest & (sgdma_tx_m_read_read);
    end


  //sgdma_tx_m_read_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_m_read_address != sgdma_tx_m_read_address_last_time))
        begin
          $write("%0d ns: sgdma_tx_m_read_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_tx_m_read_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_m_read_read_last_time <= 0;
      else 
        sgdma_tx_m_read_read_last_time <= sgdma_tx_m_read_read;
    end


  //sgdma_tx_m_read_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_m_read_read != sgdma_tx_m_read_read_last_time))
        begin
          $write("%0d ns: sgdma_tx_m_read_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_tx_out_arbitrator (
                                 // inputs:
                                  clk,
                                  reset_n,
                                  sgdma_tx_out_data,
                                  sgdma_tx_out_empty,
                                  sgdma_tx_out_endofpacket,
                                  sgdma_tx_out_error,
                                  sgdma_tx_out_startofpacket,
                                  sgdma_tx_out_valid,
                                  tse_mac_transmit_ready_from_sa,

                                 // outputs:
                                  sgdma_tx_out_ready
                               )
;

  output           sgdma_tx_out_ready;
  input            clk;
  input            reset_n;
  input   [ 31: 0] sgdma_tx_out_data;
  input   [  1: 0] sgdma_tx_out_empty;
  input            sgdma_tx_out_endofpacket;
  input            sgdma_tx_out_error;
  input            sgdma_tx_out_startofpacket;
  input            sgdma_tx_out_valid;
  input            tse_mac_transmit_ready_from_sa;

  wire             sgdma_tx_out_ready;
  //mux sgdma_tx_out_ready, which is an e_mux
  assign sgdma_tx_out_ready = tse_mac_transmit_ready_from_sa;


endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sysid_control_slave_arbitrator (
                                        // inputs:
                                         clk,
                                         pb_cpu_to_io_m1_address_to_slave,
                                         pb_cpu_to_io_m1_burstcount,
                                         pb_cpu_to_io_m1_chipselect,
                                         pb_cpu_to_io_m1_latency_counter,
                                         pb_cpu_to_io_m1_read,
                                         pb_cpu_to_io_m1_write,
                                         reset_n,
                                         sysid_control_slave_readdata,

                                        // outputs:
                                         d1_sysid_control_slave_end_xfer,
                                         pb_cpu_to_io_m1_granted_sysid_control_slave,
                                         pb_cpu_to_io_m1_qualified_request_sysid_control_slave,
                                         pb_cpu_to_io_m1_read_data_valid_sysid_control_slave,
                                         pb_cpu_to_io_m1_requests_sysid_control_slave,
                                         sysid_control_slave_address,
                                         sysid_control_slave_readdata_from_sa,
                                         sysid_control_slave_reset_n
                                      )
;

  output           d1_sysid_control_slave_end_xfer;
  output           pb_cpu_to_io_m1_granted_sysid_control_slave;
  output           pb_cpu_to_io_m1_qualified_request_sysid_control_slave;
  output           pb_cpu_to_io_m1_read_data_valid_sysid_control_slave;
  output           pb_cpu_to_io_m1_requests_sysid_control_slave;
  output           sysid_control_slave_address;
  output  [ 31: 0] sysid_control_slave_readdata_from_sa;
  output           sysid_control_slave_reset_n;
  input            clk;
  input   [ 22: 0] pb_cpu_to_io_m1_address_to_slave;
  input            pb_cpu_to_io_m1_burstcount;
  input            pb_cpu_to_io_m1_chipselect;
  input            pb_cpu_to_io_m1_latency_counter;
  input            pb_cpu_to_io_m1_read;
  input            pb_cpu_to_io_m1_write;
  input            reset_n;
  input   [ 31: 0] sysid_control_slave_readdata;

  reg              d1_reasons_to_wait;
  reg              d1_sysid_control_slave_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sysid_control_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             pb_cpu_to_io_m1_arbiterlock;
  wire             pb_cpu_to_io_m1_arbiterlock2;
  wire             pb_cpu_to_io_m1_continuerequest;
  wire             pb_cpu_to_io_m1_granted_sysid_control_slave;
  wire             pb_cpu_to_io_m1_qualified_request_sysid_control_slave;
  wire             pb_cpu_to_io_m1_read_data_valid_sysid_control_slave;
  wire             pb_cpu_to_io_m1_requests_sysid_control_slave;
  wire             pb_cpu_to_io_m1_saved_grant_sysid_control_slave;
  wire    [ 22: 0] shifted_address_to_sysid_control_slave_from_pb_cpu_to_io_m1;
  wire             sysid_control_slave_address;
  wire             sysid_control_slave_allgrants;
  wire             sysid_control_slave_allow_new_arb_cycle;
  wire             sysid_control_slave_any_bursting_master_saved_grant;
  wire             sysid_control_slave_any_continuerequest;
  wire             sysid_control_slave_arb_counter_enable;
  reg              sysid_control_slave_arb_share_counter;
  wire             sysid_control_slave_arb_share_counter_next_value;
  wire             sysid_control_slave_arb_share_set_values;
  wire             sysid_control_slave_beginbursttransfer_internal;
  wire             sysid_control_slave_begins_xfer;
  wire             sysid_control_slave_end_xfer;
  wire             sysid_control_slave_firsttransfer;
  wire             sysid_control_slave_grant_vector;
  wire             sysid_control_slave_in_a_read_cycle;
  wire             sysid_control_slave_in_a_write_cycle;
  wire             sysid_control_slave_master_qreq_vector;
  wire             sysid_control_slave_non_bursting_master_requests;
  wire    [ 31: 0] sysid_control_slave_readdata_from_sa;
  reg              sysid_control_slave_reg_firsttransfer;
  wire             sysid_control_slave_reset_n;
  reg              sysid_control_slave_slavearbiterlockenable;
  wire             sysid_control_slave_slavearbiterlockenable2;
  wire             sysid_control_slave_unreg_firsttransfer;
  wire             sysid_control_slave_waits_for_read;
  wire             sysid_control_slave_waits_for_write;
  wire             wait_for_sysid_control_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sysid_control_slave_end_xfer;
    end


  assign sysid_control_slave_begins_xfer = ~d1_reasons_to_wait & ((pb_cpu_to_io_m1_qualified_request_sysid_control_slave));
  //assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata;

  assign pb_cpu_to_io_m1_requests_sysid_control_slave = (({pb_cpu_to_io_m1_address_to_slave[22 : 3] , 3'b0} == 23'h4d40) & pb_cpu_to_io_m1_chipselect) & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect);
  //sysid_control_slave_arb_share_counter set values, which is an e_mux
  assign sysid_control_slave_arb_share_set_values = 1;

  //sysid_control_slave_non_bursting_master_requests mux, which is an e_mux
  assign sysid_control_slave_non_bursting_master_requests = pb_cpu_to_io_m1_requests_sysid_control_slave;

  //sysid_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign sysid_control_slave_any_bursting_master_saved_grant = 0;

  //sysid_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign sysid_control_slave_arb_share_counter_next_value = sysid_control_slave_firsttransfer ? (sysid_control_slave_arb_share_set_values - 1) : |sysid_control_slave_arb_share_counter ? (sysid_control_slave_arb_share_counter - 1) : 0;

  //sysid_control_slave_allgrants all slave grants, which is an e_mux
  assign sysid_control_slave_allgrants = |sysid_control_slave_grant_vector;

  //sysid_control_slave_end_xfer assignment, which is an e_assign
  assign sysid_control_slave_end_xfer = ~(sysid_control_slave_waits_for_read | sysid_control_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_sysid_control_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sysid_control_slave = sysid_control_slave_end_xfer & (~sysid_control_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sysid_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign sysid_control_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_sysid_control_slave & sysid_control_slave_allgrants) | (end_xfer_arb_share_counter_term_sysid_control_slave & ~sysid_control_slave_non_bursting_master_requests);

  //sysid_control_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_arb_share_counter <= 0;
      else if (sysid_control_slave_arb_counter_enable)
          sysid_control_slave_arb_share_counter <= sysid_control_slave_arb_share_counter_next_value;
    end


  //sysid_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_slavearbiterlockenable <= 0;
      else if ((|sysid_control_slave_master_qreq_vector & end_xfer_arb_share_counter_term_sysid_control_slave) | (end_xfer_arb_share_counter_term_sysid_control_slave & ~sysid_control_slave_non_bursting_master_requests))
          sysid_control_slave_slavearbiterlockenable <= |sysid_control_slave_arb_share_counter_next_value;
    end


  //pb_cpu_to_io/m1 sysid/control_slave arbiterlock, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock = sysid_control_slave_slavearbiterlockenable & pb_cpu_to_io_m1_continuerequest;

  //sysid_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sysid_control_slave_slavearbiterlockenable2 = |sysid_control_slave_arb_share_counter_next_value;

  //pb_cpu_to_io/m1 sysid/control_slave arbiterlock2, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock2 = sysid_control_slave_slavearbiterlockenable2 & pb_cpu_to_io_m1_continuerequest;

  //sysid_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign sysid_control_slave_any_continuerequest = 1;

  //pb_cpu_to_io_m1_continuerequest continued request, which is an e_assign
  assign pb_cpu_to_io_m1_continuerequest = 1;

  assign pb_cpu_to_io_m1_qualified_request_sysid_control_slave = pb_cpu_to_io_m1_requests_sysid_control_slave & ~(((pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ((pb_cpu_to_io_m1_latency_counter != 0))));
  //local readdatavalid pb_cpu_to_io_m1_read_data_valid_sysid_control_slave, which is an e_mux
  assign pb_cpu_to_io_m1_read_data_valid_sysid_control_slave = pb_cpu_to_io_m1_granted_sysid_control_slave & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ~sysid_control_slave_waits_for_read;

  //master is always granted when requested
  assign pb_cpu_to_io_m1_granted_sysid_control_slave = pb_cpu_to_io_m1_qualified_request_sysid_control_slave;

  //pb_cpu_to_io/m1 saved-grant sysid/control_slave, which is an e_assign
  assign pb_cpu_to_io_m1_saved_grant_sysid_control_slave = pb_cpu_to_io_m1_requests_sysid_control_slave;

  //allow new arb cycle for sysid/control_slave, which is an e_assign
  assign sysid_control_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign sysid_control_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign sysid_control_slave_master_qreq_vector = 1;

  //sysid_control_slave_reset_n assignment, which is an e_assign
  assign sysid_control_slave_reset_n = reset_n;

  //sysid_control_slave_firsttransfer first transaction, which is an e_assign
  assign sysid_control_slave_firsttransfer = sysid_control_slave_begins_xfer ? sysid_control_slave_unreg_firsttransfer : sysid_control_slave_reg_firsttransfer;

  //sysid_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign sysid_control_slave_unreg_firsttransfer = ~(sysid_control_slave_slavearbiterlockenable & sysid_control_slave_any_continuerequest);

  //sysid_control_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_reg_firsttransfer <= 1'b1;
      else if (sysid_control_slave_begins_xfer)
          sysid_control_slave_reg_firsttransfer <= sysid_control_slave_unreg_firsttransfer;
    end


  //sysid_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sysid_control_slave_beginbursttransfer_internal = sysid_control_slave_begins_xfer;

  assign shifted_address_to_sysid_control_slave_from_pb_cpu_to_io_m1 = pb_cpu_to_io_m1_address_to_slave;
  //sysid_control_slave_address mux, which is an e_mux
  assign sysid_control_slave_address = shifted_address_to_sysid_control_slave_from_pb_cpu_to_io_m1 >> 2;

  //d1_sysid_control_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sysid_control_slave_end_xfer <= 1;
      else 
        d1_sysid_control_slave_end_xfer <= sysid_control_slave_end_xfer;
    end


  //sysid_control_slave_waits_for_read in a cycle, which is an e_mux
  assign sysid_control_slave_waits_for_read = sysid_control_slave_in_a_read_cycle & sysid_control_slave_begins_xfer;

  //sysid_control_slave_in_a_read_cycle assignment, which is an e_assign
  assign sysid_control_slave_in_a_read_cycle = pb_cpu_to_io_m1_granted_sysid_control_slave & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sysid_control_slave_in_a_read_cycle;

  //sysid_control_slave_waits_for_write in a cycle, which is an e_mux
  assign sysid_control_slave_waits_for_write = sysid_control_slave_in_a_write_cycle & 0;

  //sysid_control_slave_in_a_write_cycle assignment, which is an e_assign
  assign sysid_control_slave_in_a_write_cycle = pb_cpu_to_io_m1_granted_sysid_control_slave & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sysid_control_slave_in_a_write_cycle;

  assign wait_for_sysid_control_slave_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sysid/control_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pb_cpu_to_io/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_io_m1_requests_sysid_control_slave && (pb_cpu_to_io_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pb_cpu_to_io/m1 drove 0 on its 'burstcount' port while accessing slave sysid/control_slave", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tb_fsm_avalon_slave_arbitrator (
                                        // inputs:
                                         clk,
                                         pb_cpu_to_fsm_m1_address_to_slave,
                                         pb_cpu_to_fsm_m1_burstcount,
                                         pb_cpu_to_fsm_m1_byteenable,
                                         pb_cpu_to_fsm_m1_chipselect,
                                         pb_cpu_to_fsm_m1_dbs_address,
                                         pb_cpu_to_fsm_m1_dbs_write_16,
                                         pb_cpu_to_fsm_m1_latency_counter,
                                         pb_cpu_to_fsm_m1_read,
                                         pb_cpu_to_fsm_m1_write,
                                         reset_n,

                                        // outputs:
                                         d1_tb_fsm_avalon_slave_end_xfer,
                                         ext_flash_1_s1_wait_counter_eq_0,
                                         ext_flash_s1_wait_counter_eq_0,
                                         incoming_tb_fsm_data_with_Xs_converted_to_0,
                                         pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1,
                                         pb_cpu_to_fsm_m1_byteenable_ext_flash_s1,
                                         pb_cpu_to_fsm_m1_granted_ext_flash_1_s1,
                                         pb_cpu_to_fsm_m1_granted_ext_flash_s1,
                                         pb_cpu_to_fsm_m1_qualified_request_ext_flash_1_s1,
                                         pb_cpu_to_fsm_m1_qualified_request_ext_flash_s1,
                                         pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1,
                                         pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1,
                                         pb_cpu_to_fsm_m1_requests_ext_flash_1_s1,
                                         pb_cpu_to_fsm_m1_requests_ext_flash_s1,
                                         select_n_to_the_ext_flash,
                                         select_n_to_the_ext_flash_1,
                                         tb_fsm_address,
                                         tb_fsm_data,
                                         tb_fsm_readn,
                                         tb_fsm_writen
                                      )
;

  output           d1_tb_fsm_avalon_slave_end_xfer;
  output           ext_flash_1_s1_wait_counter_eq_0;
  output           ext_flash_s1_wait_counter_eq_0;
  output  [ 15: 0] incoming_tb_fsm_data_with_Xs_converted_to_0;
  output  [  1: 0] pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1;
  output  [  1: 0] pb_cpu_to_fsm_m1_byteenable_ext_flash_s1;
  output           pb_cpu_to_fsm_m1_granted_ext_flash_1_s1;
  output           pb_cpu_to_fsm_m1_granted_ext_flash_s1;
  output           pb_cpu_to_fsm_m1_qualified_request_ext_flash_1_s1;
  output           pb_cpu_to_fsm_m1_qualified_request_ext_flash_s1;
  output           pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1;
  output           pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1;
  output           pb_cpu_to_fsm_m1_requests_ext_flash_1_s1;
  output           pb_cpu_to_fsm_m1_requests_ext_flash_s1;
  output           select_n_to_the_ext_flash;
  output           select_n_to_the_ext_flash_1;
  output  [ 24: 0] tb_fsm_address;
  inout   [ 15: 0] tb_fsm_data;
  output           tb_fsm_readn;
  output           tb_fsm_writen;
  input            clk;
  input   [ 25: 0] pb_cpu_to_fsm_m1_address_to_slave;
  input            pb_cpu_to_fsm_m1_burstcount;
  input   [  3: 0] pb_cpu_to_fsm_m1_byteenable;
  input            pb_cpu_to_fsm_m1_chipselect;
  input   [  1: 0] pb_cpu_to_fsm_m1_dbs_address;
  input   [ 15: 0] pb_cpu_to_fsm_m1_dbs_write_16;
  input   [  1: 0] pb_cpu_to_fsm_m1_latency_counter;
  input            pb_cpu_to_fsm_m1_read;
  input            pb_cpu_to_fsm_m1_write;
  input            reset_n;

  reg              d1_in_a_write_cycle /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_ENABLE_REGISTER=ON"  */;
  reg     [ 15: 0] d1_outgoing_tb_fsm_data /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              d1_reasons_to_wait;
  reg              d1_tb_fsm_avalon_slave_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_tb_fsm_avalon_slave;
  wire    [  4: 0] ext_flash_1_s1_counter_load_value;
  wire             ext_flash_1_s1_in_a_read_cycle;
  wire             ext_flash_1_s1_in_a_write_cycle;
  reg     [  4: 0] ext_flash_1_s1_wait_counter;
  wire             ext_flash_1_s1_wait_counter_eq_0;
  wire             ext_flash_1_s1_waits_for_read;
  wire             ext_flash_1_s1_waits_for_write;
  wire             ext_flash_1_s1_with_write_latency;
  wire    [  4: 0] ext_flash_s1_counter_load_value;
  wire             ext_flash_s1_in_a_read_cycle;
  wire             ext_flash_s1_in_a_write_cycle;
  reg     [  4: 0] ext_flash_s1_wait_counter;
  wire             ext_flash_s1_wait_counter_eq_0;
  wire             ext_flash_s1_waits_for_read;
  wire             ext_flash_s1_waits_for_write;
  wire             ext_flash_s1_with_write_latency;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg     [ 15: 0] incoming_tb_fsm_data /* synthesis ALTERA_ATTRIBUTE = "FAST_INPUT_REGISTER=ON"  */;
  wire             incoming_tb_fsm_data_bit_0_is_x;
  wire             incoming_tb_fsm_data_bit_10_is_x;
  wire             incoming_tb_fsm_data_bit_11_is_x;
  wire             incoming_tb_fsm_data_bit_12_is_x;
  wire             incoming_tb_fsm_data_bit_13_is_x;
  wire             incoming_tb_fsm_data_bit_14_is_x;
  wire             incoming_tb_fsm_data_bit_15_is_x;
  wire             incoming_tb_fsm_data_bit_1_is_x;
  wire             incoming_tb_fsm_data_bit_2_is_x;
  wire             incoming_tb_fsm_data_bit_3_is_x;
  wire             incoming_tb_fsm_data_bit_4_is_x;
  wire             incoming_tb_fsm_data_bit_5_is_x;
  wire             incoming_tb_fsm_data_bit_6_is_x;
  wire             incoming_tb_fsm_data_bit_7_is_x;
  wire             incoming_tb_fsm_data_bit_8_is_x;
  wire             incoming_tb_fsm_data_bit_9_is_x;
  wire    [ 15: 0] incoming_tb_fsm_data_with_Xs_converted_to_0;
  wire    [ 15: 0] outgoing_tb_fsm_data;
  wire    [  1: 0] p1_pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1_shift_register;
  wire    [  1: 0] p1_pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1_shift_register;
  wire             p1_select_n_to_the_ext_flash;
  wire             p1_select_n_to_the_ext_flash_1;
  wire    [ 24: 0] p1_tb_fsm_address;
  wire             p1_tb_fsm_readn;
  wire             p1_tb_fsm_writen;
  wire             pb_cpu_to_fsm_m1_arbiterlock;
  wire             pb_cpu_to_fsm_m1_arbiterlock2;
  wire    [  1: 0] pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1;
  wire    [  1: 0] pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1_segment_0;
  wire    [  1: 0] pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1_segment_1;
  wire    [  1: 0] pb_cpu_to_fsm_m1_byteenable_ext_flash_s1;
  wire    [  1: 0] pb_cpu_to_fsm_m1_byteenable_ext_flash_s1_segment_0;
  wire    [  1: 0] pb_cpu_to_fsm_m1_byteenable_ext_flash_s1_segment_1;
  wire             pb_cpu_to_fsm_m1_continuerequest;
  wire             pb_cpu_to_fsm_m1_granted_ext_flash_1_s1;
  wire             pb_cpu_to_fsm_m1_granted_ext_flash_s1;
  wire             pb_cpu_to_fsm_m1_qualified_request_ext_flash_1_s1;
  wire             pb_cpu_to_fsm_m1_qualified_request_ext_flash_s1;
  wire             pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1;
  reg     [  1: 0] pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1_shift_register;
  wire             pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1_shift_register_in;
  wire             pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1;
  reg     [  1: 0] pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1_shift_register;
  wire             pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1_shift_register_in;
  wire             pb_cpu_to_fsm_m1_requests_ext_flash_1_s1;
  wire             pb_cpu_to_fsm_m1_requests_ext_flash_s1;
  wire             pb_cpu_to_fsm_m1_saved_grant_ext_flash_1_s1;
  wire             pb_cpu_to_fsm_m1_saved_grant_ext_flash_s1;
  reg              select_n_to_the_ext_flash /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              select_n_to_the_ext_flash_1 /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg     [ 24: 0] tb_fsm_address /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             tb_fsm_avalon_slave_allgrants;
  wire             tb_fsm_avalon_slave_allow_new_arb_cycle;
  wire             tb_fsm_avalon_slave_any_bursting_master_saved_grant;
  wire             tb_fsm_avalon_slave_any_continuerequest;
  wire             tb_fsm_avalon_slave_arb_counter_enable;
  reg     [  1: 0] tb_fsm_avalon_slave_arb_share_counter;
  wire    [  1: 0] tb_fsm_avalon_slave_arb_share_counter_next_value;
  wire    [  1: 0] tb_fsm_avalon_slave_arb_share_set_values;
  wire             tb_fsm_avalon_slave_beginbursttransfer_internal;
  wire             tb_fsm_avalon_slave_begins_xfer;
  wire             tb_fsm_avalon_slave_end_xfer;
  wire             tb_fsm_avalon_slave_firsttransfer;
  wire             tb_fsm_avalon_slave_grant_vector;
  wire             tb_fsm_avalon_slave_master_qreq_vector;
  wire             tb_fsm_avalon_slave_non_bursting_master_requests;
  wire             tb_fsm_avalon_slave_read_pending;
  reg              tb_fsm_avalon_slave_reg_firsttransfer;
  reg              tb_fsm_avalon_slave_slavearbiterlockenable;
  wire             tb_fsm_avalon_slave_slavearbiterlockenable2;
  wire             tb_fsm_avalon_slave_unreg_firsttransfer;
  wire             tb_fsm_avalon_slave_write_pending;
  wire    [ 15: 0] tb_fsm_data;
  reg              tb_fsm_readn /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              tb_fsm_writen /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             time_to_write;
  wire             wait_for_ext_flash_1_s1_counter;
  wire             wait_for_ext_flash_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~tb_fsm_avalon_slave_end_xfer;
    end


  assign tb_fsm_avalon_slave_begins_xfer = ~d1_reasons_to_wait & ((pb_cpu_to_fsm_m1_qualified_request_ext_flash_1_s1 | pb_cpu_to_fsm_m1_qualified_request_ext_flash_s1));
  assign pb_cpu_to_fsm_m1_requests_ext_flash_1_s1 = ({pb_cpu_to_fsm_m1_address_to_slave[25] , 25'b0} == 26'h2000000) & pb_cpu_to_fsm_m1_chipselect;
  //~select_n_to_the_ext_flash_1 of type chipselect to ~p1_select_n_to_the_ext_flash_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          select_n_to_the_ext_flash_1 <= ~0;
      else 
        select_n_to_the_ext_flash_1 <= p1_select_n_to_the_ext_flash_1;
    end


  //~select_n_to_the_ext_flash of type chipselect to ~p1_select_n_to_the_ext_flash, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          select_n_to_the_ext_flash <= ~0;
      else 
        select_n_to_the_ext_flash <= p1_select_n_to_the_ext_flash;
    end


  assign tb_fsm_avalon_slave_write_pending = 0;
  //tb_fsm/avalon_slave read pending calc, which is an e_assign
  assign tb_fsm_avalon_slave_read_pending = 0;

  //tb_fsm_avalon_slave_arb_share_counter set values, which is an e_mux
  assign tb_fsm_avalon_slave_arb_share_set_values = (pb_cpu_to_fsm_m1_granted_ext_flash_1_s1)? 2 :
    (pb_cpu_to_fsm_m1_granted_ext_flash_s1)? 2 :
    1;

  //tb_fsm_avalon_slave_non_bursting_master_requests mux, which is an e_mux
  assign tb_fsm_avalon_slave_non_bursting_master_requests = pb_cpu_to_fsm_m1_requests_ext_flash_1_s1 |
    pb_cpu_to_fsm_m1_requests_ext_flash_s1;

  //tb_fsm_avalon_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign tb_fsm_avalon_slave_any_bursting_master_saved_grant = 0;

  //tb_fsm_avalon_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign tb_fsm_avalon_slave_arb_share_counter_next_value = tb_fsm_avalon_slave_firsttransfer ? (tb_fsm_avalon_slave_arb_share_set_values - 1) : |tb_fsm_avalon_slave_arb_share_counter ? (tb_fsm_avalon_slave_arb_share_counter - 1) : 0;

  //tb_fsm_avalon_slave_allgrants all slave grants, which is an e_mux
  assign tb_fsm_avalon_slave_allgrants = (|tb_fsm_avalon_slave_grant_vector) |
    (|tb_fsm_avalon_slave_grant_vector);

  //tb_fsm_avalon_slave_end_xfer assignment, which is an e_assign
  assign tb_fsm_avalon_slave_end_xfer = ~(ext_flash_1_s1_waits_for_read | ext_flash_1_s1_waits_for_write | ext_flash_s1_waits_for_read | ext_flash_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_tb_fsm_avalon_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_tb_fsm_avalon_slave = tb_fsm_avalon_slave_end_xfer & (~tb_fsm_avalon_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //tb_fsm_avalon_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign tb_fsm_avalon_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_tb_fsm_avalon_slave & tb_fsm_avalon_slave_allgrants) | (end_xfer_arb_share_counter_term_tb_fsm_avalon_slave & ~tb_fsm_avalon_slave_non_bursting_master_requests);

  //tb_fsm_avalon_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tb_fsm_avalon_slave_arb_share_counter <= 0;
      else if (tb_fsm_avalon_slave_arb_counter_enable)
          tb_fsm_avalon_slave_arb_share_counter <= tb_fsm_avalon_slave_arb_share_counter_next_value;
    end


  //tb_fsm_avalon_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tb_fsm_avalon_slave_slavearbiterlockenable <= 0;
      else if ((|tb_fsm_avalon_slave_master_qreq_vector & end_xfer_arb_share_counter_term_tb_fsm_avalon_slave) | (end_xfer_arb_share_counter_term_tb_fsm_avalon_slave & ~tb_fsm_avalon_slave_non_bursting_master_requests))
          tb_fsm_avalon_slave_slavearbiterlockenable <= |tb_fsm_avalon_slave_arb_share_counter_next_value;
    end


  //pb_cpu_to_fsm/m1 tb_fsm/avalon_slave arbiterlock, which is an e_assign
  assign pb_cpu_to_fsm_m1_arbiterlock = tb_fsm_avalon_slave_slavearbiterlockenable & pb_cpu_to_fsm_m1_continuerequest;

  //tb_fsm_avalon_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign tb_fsm_avalon_slave_slavearbiterlockenable2 = |tb_fsm_avalon_slave_arb_share_counter_next_value;

  //pb_cpu_to_fsm/m1 tb_fsm/avalon_slave arbiterlock2, which is an e_assign
  assign pb_cpu_to_fsm_m1_arbiterlock2 = tb_fsm_avalon_slave_slavearbiterlockenable2 & pb_cpu_to_fsm_m1_continuerequest;

  //tb_fsm_avalon_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign tb_fsm_avalon_slave_any_continuerequest = 1;

  //pb_cpu_to_fsm_m1_continuerequest continued request, which is an e_assign
  assign pb_cpu_to_fsm_m1_continuerequest = 1;

  assign pb_cpu_to_fsm_m1_qualified_request_ext_flash_1_s1 = pb_cpu_to_fsm_m1_requests_ext_flash_1_s1 & ~(((pb_cpu_to_fsm_m1_read & pb_cpu_to_fsm_m1_chipselect) & (tb_fsm_avalon_slave_write_pending | (tb_fsm_avalon_slave_read_pending) | (2 < pb_cpu_to_fsm_m1_latency_counter))) | ((tb_fsm_avalon_slave_read_pending | !pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1) & (pb_cpu_to_fsm_m1_write & pb_cpu_to_fsm_m1_chipselect)));
  //pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1_shift_register_in = pb_cpu_to_fsm_m1_granted_ext_flash_1_s1 & (pb_cpu_to_fsm_m1_read & pb_cpu_to_fsm_m1_chipselect) & ~ext_flash_1_s1_waits_for_read;

  //shift register p1 pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1_shift_register = {pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1_shift_register, pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1_shift_register_in};

  //pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1_shift_register <= 0;
      else 
        pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1_shift_register <= p1_pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1_shift_register;
    end


  //local readdatavalid pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1, which is an e_mux
  assign pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1 = pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1_shift_register[1];

  //tb_fsm_data register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          incoming_tb_fsm_data <= 0;
      else 
        incoming_tb_fsm_data <= tb_fsm_data;
    end


  //ext_flash_1_s1_with_write_latency assignment, which is an e_assign
  assign ext_flash_1_s1_with_write_latency = in_a_write_cycle & (pb_cpu_to_fsm_m1_qualified_request_ext_flash_1_s1);

  //time to write the data, which is an e_mux
  assign time_to_write = (ext_flash_1_s1_with_write_latency)? 1 :
    (ext_flash_s1_with_write_latency)? 1 :
    0;

  //d1_outgoing_tb_fsm_data register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_outgoing_tb_fsm_data <= 0;
      else 
        d1_outgoing_tb_fsm_data <= outgoing_tb_fsm_data;
    end


  //write cycle delayed by 1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_in_a_write_cycle <= 0;
      else 
        d1_in_a_write_cycle <= time_to_write;
    end


  //d1_outgoing_tb_fsm_data tristate driver, which is an e_assign
  assign tb_fsm_data = (d1_in_a_write_cycle)? d1_outgoing_tb_fsm_data:{16{1'bz}};

  //outgoing_tb_fsm_data mux, which is an e_mux
  assign outgoing_tb_fsm_data = (pb_cpu_to_fsm_m1_granted_ext_flash_1_s1)? pb_cpu_to_fsm_m1_dbs_write_16 :
    pb_cpu_to_fsm_m1_dbs_write_16;

  assign pb_cpu_to_fsm_m1_requests_ext_flash_s1 = ({pb_cpu_to_fsm_m1_address_to_slave[25] , 25'b0} == 26'h0) & pb_cpu_to_fsm_m1_chipselect;
  assign pb_cpu_to_fsm_m1_qualified_request_ext_flash_s1 = pb_cpu_to_fsm_m1_requests_ext_flash_s1 & ~(((pb_cpu_to_fsm_m1_read & pb_cpu_to_fsm_m1_chipselect) & (tb_fsm_avalon_slave_write_pending | (tb_fsm_avalon_slave_read_pending) | (2 < pb_cpu_to_fsm_m1_latency_counter))) | ((tb_fsm_avalon_slave_read_pending | !pb_cpu_to_fsm_m1_byteenable_ext_flash_s1) & (pb_cpu_to_fsm_m1_write & pb_cpu_to_fsm_m1_chipselect)));
  //pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1_shift_register_in = pb_cpu_to_fsm_m1_granted_ext_flash_s1 & (pb_cpu_to_fsm_m1_read & pb_cpu_to_fsm_m1_chipselect) & ~ext_flash_s1_waits_for_read;

  //shift register p1 pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1_shift_register = {pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1_shift_register, pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1_shift_register_in};

  //pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1_shift_register <= 0;
      else 
        pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1_shift_register <= p1_pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1_shift_register;
    end


  //local readdatavalid pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1, which is an e_mux
  assign pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1 = pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1_shift_register[1];

  //ext_flash_s1_with_write_latency assignment, which is an e_assign
  assign ext_flash_s1_with_write_latency = in_a_write_cycle & (pb_cpu_to_fsm_m1_qualified_request_ext_flash_s1);

  //master is always granted when requested
  assign pb_cpu_to_fsm_m1_granted_ext_flash_1_s1 = pb_cpu_to_fsm_m1_qualified_request_ext_flash_1_s1;

  //pb_cpu_to_fsm/m1 saved-grant ext_flash_1/s1, which is an e_assign
  assign pb_cpu_to_fsm_m1_saved_grant_ext_flash_1_s1 = pb_cpu_to_fsm_m1_requests_ext_flash_1_s1;

  //allow new arb cycle for tb_fsm/avalon_slave, which is an e_assign
  assign tb_fsm_avalon_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign tb_fsm_avalon_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign tb_fsm_avalon_slave_master_qreq_vector = 1;

  //master is always granted when requested
  assign pb_cpu_to_fsm_m1_granted_ext_flash_s1 = pb_cpu_to_fsm_m1_qualified_request_ext_flash_s1;

  //pb_cpu_to_fsm/m1 saved-grant ext_flash/s1, which is an e_assign
  assign pb_cpu_to_fsm_m1_saved_grant_ext_flash_s1 = pb_cpu_to_fsm_m1_requests_ext_flash_s1;

  assign p1_select_n_to_the_ext_flash_1 = ~pb_cpu_to_fsm_m1_granted_ext_flash_1_s1;
  //tb_fsm_avalon_slave_firsttransfer first transaction, which is an e_assign
  assign tb_fsm_avalon_slave_firsttransfer = tb_fsm_avalon_slave_begins_xfer ? tb_fsm_avalon_slave_unreg_firsttransfer : tb_fsm_avalon_slave_reg_firsttransfer;

  //tb_fsm_avalon_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign tb_fsm_avalon_slave_unreg_firsttransfer = ~(tb_fsm_avalon_slave_slavearbiterlockenable & tb_fsm_avalon_slave_any_continuerequest);

  //tb_fsm_avalon_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tb_fsm_avalon_slave_reg_firsttransfer <= 1'b1;
      else if (tb_fsm_avalon_slave_begins_xfer)
          tb_fsm_avalon_slave_reg_firsttransfer <= tb_fsm_avalon_slave_unreg_firsttransfer;
    end


  //tb_fsm_avalon_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign tb_fsm_avalon_slave_beginbursttransfer_internal = tb_fsm_avalon_slave_begins_xfer;

  //~tb_fsm_readn of type read to ~p1_tb_fsm_readn, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tb_fsm_readn <= ~0;
      else 
        tb_fsm_readn <= p1_tb_fsm_readn;
    end


  //~p1_tb_fsm_readn assignment, which is an e_mux
  assign p1_tb_fsm_readn = ~((((pb_cpu_to_fsm_m1_granted_ext_flash_1_s1 & (pb_cpu_to_fsm_m1_read & pb_cpu_to_fsm_m1_chipselect)))& ~tb_fsm_avalon_slave_begins_xfer & (ext_flash_1_s1_wait_counter < 16)) |
    (((pb_cpu_to_fsm_m1_granted_ext_flash_s1 & (pb_cpu_to_fsm_m1_read & pb_cpu_to_fsm_m1_chipselect)))& ~tb_fsm_avalon_slave_begins_xfer & (ext_flash_s1_wait_counter < 16)));

  //~tb_fsm_writen of type write to ~p1_tb_fsm_writen, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tb_fsm_writen <= ~0;
      else 
        tb_fsm_writen <= p1_tb_fsm_writen;
    end


  //~p1_tb_fsm_writen assignment, which is an e_mux
  assign p1_tb_fsm_writen = ~(((((pb_cpu_to_fsm_m1_granted_ext_flash_1_s1 & (pb_cpu_to_fsm_m1_write & pb_cpu_to_fsm_m1_chipselect))) & ~tb_fsm_avalon_slave_begins_xfer & (ext_flash_1_s1_wait_counter >= 3) & (ext_flash_1_s1_wait_counter < 19))) |
    ((((pb_cpu_to_fsm_m1_granted_ext_flash_s1 & (pb_cpu_to_fsm_m1_write & pb_cpu_to_fsm_m1_chipselect))) & ~tb_fsm_avalon_slave_begins_xfer & (ext_flash_s1_wait_counter >= 3) & (ext_flash_s1_wait_counter < 19))));

  //tb_fsm_address of type address to p1_tb_fsm_address, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tb_fsm_address <= 0;
      else 
        tb_fsm_address <= p1_tb_fsm_address;
    end


  //p1_tb_fsm_address mux, which is an e_mux
  assign p1_tb_fsm_address = (pb_cpu_to_fsm_m1_granted_ext_flash_1_s1)? ({pb_cpu_to_fsm_m1_address_to_slave >> 2,
    pb_cpu_to_fsm_m1_dbs_address[1],
    {1 {1'b0}}}) :
    ({pb_cpu_to_fsm_m1_address_to_slave >> 2,
    pb_cpu_to_fsm_m1_dbs_address[1],
    {1 {1'b0}}});

  //d1_tb_fsm_avalon_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_tb_fsm_avalon_slave_end_xfer <= 1;
      else 
        d1_tb_fsm_avalon_slave_end_xfer <= tb_fsm_avalon_slave_end_xfer;
    end


  //ext_flash_1_s1_waits_for_read in a cycle, which is an e_mux
  assign ext_flash_1_s1_waits_for_read = ext_flash_1_s1_in_a_read_cycle & wait_for_ext_flash_1_s1_counter;

  //ext_flash_1_s1_in_a_read_cycle assignment, which is an e_assign
  assign ext_flash_1_s1_in_a_read_cycle = pb_cpu_to_fsm_m1_granted_ext_flash_1_s1 & (pb_cpu_to_fsm_m1_read & pb_cpu_to_fsm_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = ext_flash_1_s1_in_a_read_cycle |
    ext_flash_s1_in_a_read_cycle;

  //ext_flash_1_s1_waits_for_write in a cycle, which is an e_mux
  assign ext_flash_1_s1_waits_for_write = ext_flash_1_s1_in_a_write_cycle & wait_for_ext_flash_1_s1_counter;

  //ext_flash_1_s1_in_a_write_cycle assignment, which is an e_assign
  assign ext_flash_1_s1_in_a_write_cycle = pb_cpu_to_fsm_m1_granted_ext_flash_1_s1 & (pb_cpu_to_fsm_m1_write & pb_cpu_to_fsm_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = ext_flash_1_s1_in_a_write_cycle |
    ext_flash_s1_in_a_write_cycle;

  assign ext_flash_1_s1_wait_counter_eq_0 = ext_flash_1_s1_wait_counter == 0;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_flash_1_s1_wait_counter <= 0;
      else 
        ext_flash_1_s1_wait_counter <= ext_flash_1_s1_counter_load_value;
    end


  assign ext_flash_1_s1_counter_load_value = ((ext_flash_1_s1_in_a_read_cycle & tb_fsm_avalon_slave_begins_xfer))? 18 :
    ((ext_flash_1_s1_in_a_write_cycle & tb_fsm_avalon_slave_begins_xfer))? 21 :
    (~ext_flash_1_s1_wait_counter_eq_0)? ext_flash_1_s1_wait_counter - 1 :
    0;

  assign wait_for_ext_flash_1_s1_counter = tb_fsm_avalon_slave_begins_xfer | ~ext_flash_1_s1_wait_counter_eq_0;
  assign {pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1_segment_1,
pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1_segment_0} = pb_cpu_to_fsm_m1_byteenable;
  assign pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1 = ((pb_cpu_to_fsm_m1_dbs_address[1] == 0))? pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1_segment_0 :
    pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1_segment_1;

  assign p1_select_n_to_the_ext_flash = ~pb_cpu_to_fsm_m1_granted_ext_flash_s1;
  //ext_flash_s1_waits_for_read in a cycle, which is an e_mux
  assign ext_flash_s1_waits_for_read = ext_flash_s1_in_a_read_cycle & wait_for_ext_flash_s1_counter;

  //ext_flash_s1_in_a_read_cycle assignment, which is an e_assign
  assign ext_flash_s1_in_a_read_cycle = pb_cpu_to_fsm_m1_granted_ext_flash_s1 & (pb_cpu_to_fsm_m1_read & pb_cpu_to_fsm_m1_chipselect);

  //ext_flash_s1_waits_for_write in a cycle, which is an e_mux
  assign ext_flash_s1_waits_for_write = ext_flash_s1_in_a_write_cycle & wait_for_ext_flash_s1_counter;

  //ext_flash_s1_in_a_write_cycle assignment, which is an e_assign
  assign ext_flash_s1_in_a_write_cycle = pb_cpu_to_fsm_m1_granted_ext_flash_s1 & (pb_cpu_to_fsm_m1_write & pb_cpu_to_fsm_m1_chipselect);

  assign ext_flash_s1_wait_counter_eq_0 = ext_flash_s1_wait_counter == 0;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_flash_s1_wait_counter <= 0;
      else 
        ext_flash_s1_wait_counter <= ext_flash_s1_counter_load_value;
    end


  assign ext_flash_s1_counter_load_value = ((ext_flash_s1_in_a_read_cycle & tb_fsm_avalon_slave_begins_xfer))? 18 :
    ((ext_flash_s1_in_a_write_cycle & tb_fsm_avalon_slave_begins_xfer))? 21 :
    (~ext_flash_s1_wait_counter_eq_0)? ext_flash_s1_wait_counter - 1 :
    0;

  assign wait_for_ext_flash_s1_counter = tb_fsm_avalon_slave_begins_xfer | ~ext_flash_s1_wait_counter_eq_0;
  assign {pb_cpu_to_fsm_m1_byteenable_ext_flash_s1_segment_1,
pb_cpu_to_fsm_m1_byteenable_ext_flash_s1_segment_0} = pb_cpu_to_fsm_m1_byteenable;
  assign pb_cpu_to_fsm_m1_byteenable_ext_flash_s1 = ((pb_cpu_to_fsm_m1_dbs_address[1] == 0))? pb_cpu_to_fsm_m1_byteenable_ext_flash_s1_segment_0 :
    pb_cpu_to_fsm_m1_byteenable_ext_flash_s1_segment_1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //incoming_tb_fsm_data_bit_0_is_x x check, which is an e_assign_is_x
  assign incoming_tb_fsm_data_bit_0_is_x = ^(incoming_tb_fsm_data[0]) === 1'bx;

  //Crush incoming_tb_fsm_data_with_Xs_converted_to_0[0] Xs to 0, which is an e_assign
  assign incoming_tb_fsm_data_with_Xs_converted_to_0[0] = incoming_tb_fsm_data_bit_0_is_x ? 1'b0 : incoming_tb_fsm_data[0];

  //incoming_tb_fsm_data_bit_1_is_x x check, which is an e_assign_is_x
  assign incoming_tb_fsm_data_bit_1_is_x = ^(incoming_tb_fsm_data[1]) === 1'bx;

  //Crush incoming_tb_fsm_data_with_Xs_converted_to_0[1] Xs to 0, which is an e_assign
  assign incoming_tb_fsm_data_with_Xs_converted_to_0[1] = incoming_tb_fsm_data_bit_1_is_x ? 1'b0 : incoming_tb_fsm_data[1];

  //incoming_tb_fsm_data_bit_2_is_x x check, which is an e_assign_is_x
  assign incoming_tb_fsm_data_bit_2_is_x = ^(incoming_tb_fsm_data[2]) === 1'bx;

  //Crush incoming_tb_fsm_data_with_Xs_converted_to_0[2] Xs to 0, which is an e_assign
  assign incoming_tb_fsm_data_with_Xs_converted_to_0[2] = incoming_tb_fsm_data_bit_2_is_x ? 1'b0 : incoming_tb_fsm_data[2];

  //incoming_tb_fsm_data_bit_3_is_x x check, which is an e_assign_is_x
  assign incoming_tb_fsm_data_bit_3_is_x = ^(incoming_tb_fsm_data[3]) === 1'bx;

  //Crush incoming_tb_fsm_data_with_Xs_converted_to_0[3] Xs to 0, which is an e_assign
  assign incoming_tb_fsm_data_with_Xs_converted_to_0[3] = incoming_tb_fsm_data_bit_3_is_x ? 1'b0 : incoming_tb_fsm_data[3];

  //incoming_tb_fsm_data_bit_4_is_x x check, which is an e_assign_is_x
  assign incoming_tb_fsm_data_bit_4_is_x = ^(incoming_tb_fsm_data[4]) === 1'bx;

  //Crush incoming_tb_fsm_data_with_Xs_converted_to_0[4] Xs to 0, which is an e_assign
  assign incoming_tb_fsm_data_with_Xs_converted_to_0[4] = incoming_tb_fsm_data_bit_4_is_x ? 1'b0 : incoming_tb_fsm_data[4];

  //incoming_tb_fsm_data_bit_5_is_x x check, which is an e_assign_is_x
  assign incoming_tb_fsm_data_bit_5_is_x = ^(incoming_tb_fsm_data[5]) === 1'bx;

  //Crush incoming_tb_fsm_data_with_Xs_converted_to_0[5] Xs to 0, which is an e_assign
  assign incoming_tb_fsm_data_with_Xs_converted_to_0[5] = incoming_tb_fsm_data_bit_5_is_x ? 1'b0 : incoming_tb_fsm_data[5];

  //incoming_tb_fsm_data_bit_6_is_x x check, which is an e_assign_is_x
  assign incoming_tb_fsm_data_bit_6_is_x = ^(incoming_tb_fsm_data[6]) === 1'bx;

  //Crush incoming_tb_fsm_data_with_Xs_converted_to_0[6] Xs to 0, which is an e_assign
  assign incoming_tb_fsm_data_with_Xs_converted_to_0[6] = incoming_tb_fsm_data_bit_6_is_x ? 1'b0 : incoming_tb_fsm_data[6];

  //incoming_tb_fsm_data_bit_7_is_x x check, which is an e_assign_is_x
  assign incoming_tb_fsm_data_bit_7_is_x = ^(incoming_tb_fsm_data[7]) === 1'bx;

  //Crush incoming_tb_fsm_data_with_Xs_converted_to_0[7] Xs to 0, which is an e_assign
  assign incoming_tb_fsm_data_with_Xs_converted_to_0[7] = incoming_tb_fsm_data_bit_7_is_x ? 1'b0 : incoming_tb_fsm_data[7];

  //incoming_tb_fsm_data_bit_8_is_x x check, which is an e_assign_is_x
  assign incoming_tb_fsm_data_bit_8_is_x = ^(incoming_tb_fsm_data[8]) === 1'bx;

  //Crush incoming_tb_fsm_data_with_Xs_converted_to_0[8] Xs to 0, which is an e_assign
  assign incoming_tb_fsm_data_with_Xs_converted_to_0[8] = incoming_tb_fsm_data_bit_8_is_x ? 1'b0 : incoming_tb_fsm_data[8];

  //incoming_tb_fsm_data_bit_9_is_x x check, which is an e_assign_is_x
  assign incoming_tb_fsm_data_bit_9_is_x = ^(incoming_tb_fsm_data[9]) === 1'bx;

  //Crush incoming_tb_fsm_data_with_Xs_converted_to_0[9] Xs to 0, which is an e_assign
  assign incoming_tb_fsm_data_with_Xs_converted_to_0[9] = incoming_tb_fsm_data_bit_9_is_x ? 1'b0 : incoming_tb_fsm_data[9];

  //incoming_tb_fsm_data_bit_10_is_x x check, which is an e_assign_is_x
  assign incoming_tb_fsm_data_bit_10_is_x = ^(incoming_tb_fsm_data[10]) === 1'bx;

  //Crush incoming_tb_fsm_data_with_Xs_converted_to_0[10] Xs to 0, which is an e_assign
  assign incoming_tb_fsm_data_with_Xs_converted_to_0[10] = incoming_tb_fsm_data_bit_10_is_x ? 1'b0 : incoming_tb_fsm_data[10];

  //incoming_tb_fsm_data_bit_11_is_x x check, which is an e_assign_is_x
  assign incoming_tb_fsm_data_bit_11_is_x = ^(incoming_tb_fsm_data[11]) === 1'bx;

  //Crush incoming_tb_fsm_data_with_Xs_converted_to_0[11] Xs to 0, which is an e_assign
  assign incoming_tb_fsm_data_with_Xs_converted_to_0[11] = incoming_tb_fsm_data_bit_11_is_x ? 1'b0 : incoming_tb_fsm_data[11];

  //incoming_tb_fsm_data_bit_12_is_x x check, which is an e_assign_is_x
  assign incoming_tb_fsm_data_bit_12_is_x = ^(incoming_tb_fsm_data[12]) === 1'bx;

  //Crush incoming_tb_fsm_data_with_Xs_converted_to_0[12] Xs to 0, which is an e_assign
  assign incoming_tb_fsm_data_with_Xs_converted_to_0[12] = incoming_tb_fsm_data_bit_12_is_x ? 1'b0 : incoming_tb_fsm_data[12];

  //incoming_tb_fsm_data_bit_13_is_x x check, which is an e_assign_is_x
  assign incoming_tb_fsm_data_bit_13_is_x = ^(incoming_tb_fsm_data[13]) === 1'bx;

  //Crush incoming_tb_fsm_data_with_Xs_converted_to_0[13] Xs to 0, which is an e_assign
  assign incoming_tb_fsm_data_with_Xs_converted_to_0[13] = incoming_tb_fsm_data_bit_13_is_x ? 1'b0 : incoming_tb_fsm_data[13];

  //incoming_tb_fsm_data_bit_14_is_x x check, which is an e_assign_is_x
  assign incoming_tb_fsm_data_bit_14_is_x = ^(incoming_tb_fsm_data[14]) === 1'bx;

  //Crush incoming_tb_fsm_data_with_Xs_converted_to_0[14] Xs to 0, which is an e_assign
  assign incoming_tb_fsm_data_with_Xs_converted_to_0[14] = incoming_tb_fsm_data_bit_14_is_x ? 1'b0 : incoming_tb_fsm_data[14];

  //incoming_tb_fsm_data_bit_15_is_x x check, which is an e_assign_is_x
  assign incoming_tb_fsm_data_bit_15_is_x = ^(incoming_tb_fsm_data[15]) === 1'bx;

  //Crush incoming_tb_fsm_data_with_Xs_converted_to_0[15] Xs to 0, which is an e_assign
  assign incoming_tb_fsm_data_with_Xs_converted_to_0[15] = incoming_tb_fsm_data_bit_15_is_x ? 1'b0 : incoming_tb_fsm_data[15];

  //ext_flash_1/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pb_cpu_to_fsm/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_fsm_m1_requests_ext_flash_1_s1 && (pb_cpu_to_fsm_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pb_cpu_to_fsm/m1 drove 0 on its 'burstcount' port while accessing slave ext_flash_1/s1", $time);
          $stop;
        end
    end


  //ext_flash/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_fsm_m1_granted_ext_flash_1_s1 + pb_cpu_to_fsm_m1_granted_ext_flash_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_fsm_m1_saved_grant_ext_flash_1_s1 + pb_cpu_to_fsm_m1_saved_grant_ext_flash_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  
//  assign incoming_tb_fsm_data_with_Xs_converted_to_0 = incoming_tb_fsm_data;
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tb_fsm_bridge_arbitrator 
;



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module timer_1ms_s1_arbitrator (
                                 // inputs:
                                  clk,
                                  pb_cpu_to_io_m1_address_to_slave,
                                  pb_cpu_to_io_m1_burstcount,
                                  pb_cpu_to_io_m1_chipselect,
                                  pb_cpu_to_io_m1_latency_counter,
                                  pb_cpu_to_io_m1_read,
                                  pb_cpu_to_io_m1_write,
                                  pb_cpu_to_io_m1_writedata,
                                  reset_n,
                                  timer_1ms_s1_irq,
                                  timer_1ms_s1_readdata,

                                 // outputs:
                                  d1_timer_1ms_s1_end_xfer,
                                  pb_cpu_to_io_m1_granted_timer_1ms_s1,
                                  pb_cpu_to_io_m1_qualified_request_timer_1ms_s1,
                                  pb_cpu_to_io_m1_read_data_valid_timer_1ms_s1,
                                  pb_cpu_to_io_m1_requests_timer_1ms_s1,
                                  timer_1ms_s1_address,
                                  timer_1ms_s1_chipselect,
                                  timer_1ms_s1_irq_from_sa,
                                  timer_1ms_s1_readdata_from_sa,
                                  timer_1ms_s1_reset_n,
                                  timer_1ms_s1_write_n,
                                  timer_1ms_s1_writedata
                               )
;

  output           d1_timer_1ms_s1_end_xfer;
  output           pb_cpu_to_io_m1_granted_timer_1ms_s1;
  output           pb_cpu_to_io_m1_qualified_request_timer_1ms_s1;
  output           pb_cpu_to_io_m1_read_data_valid_timer_1ms_s1;
  output           pb_cpu_to_io_m1_requests_timer_1ms_s1;
  output  [  2: 0] timer_1ms_s1_address;
  output           timer_1ms_s1_chipselect;
  output           timer_1ms_s1_irq_from_sa;
  output  [ 15: 0] timer_1ms_s1_readdata_from_sa;
  output           timer_1ms_s1_reset_n;
  output           timer_1ms_s1_write_n;
  output  [ 15: 0] timer_1ms_s1_writedata;
  input            clk;
  input   [ 22: 0] pb_cpu_to_io_m1_address_to_slave;
  input            pb_cpu_to_io_m1_burstcount;
  input            pb_cpu_to_io_m1_chipselect;
  input            pb_cpu_to_io_m1_latency_counter;
  input            pb_cpu_to_io_m1_read;
  input            pb_cpu_to_io_m1_write;
  input   [ 31: 0] pb_cpu_to_io_m1_writedata;
  input            reset_n;
  input            timer_1ms_s1_irq;
  input   [ 15: 0] timer_1ms_s1_readdata;

  reg              d1_reasons_to_wait;
  reg              d1_timer_1ms_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_timer_1ms_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             pb_cpu_to_io_m1_arbiterlock;
  wire             pb_cpu_to_io_m1_arbiterlock2;
  wire             pb_cpu_to_io_m1_continuerequest;
  wire             pb_cpu_to_io_m1_granted_timer_1ms_s1;
  wire             pb_cpu_to_io_m1_qualified_request_timer_1ms_s1;
  wire             pb_cpu_to_io_m1_read_data_valid_timer_1ms_s1;
  wire             pb_cpu_to_io_m1_requests_timer_1ms_s1;
  wire             pb_cpu_to_io_m1_saved_grant_timer_1ms_s1;
  wire    [ 22: 0] shifted_address_to_timer_1ms_s1_from_pb_cpu_to_io_m1;
  wire    [  2: 0] timer_1ms_s1_address;
  wire             timer_1ms_s1_allgrants;
  wire             timer_1ms_s1_allow_new_arb_cycle;
  wire             timer_1ms_s1_any_bursting_master_saved_grant;
  wire             timer_1ms_s1_any_continuerequest;
  wire             timer_1ms_s1_arb_counter_enable;
  reg              timer_1ms_s1_arb_share_counter;
  wire             timer_1ms_s1_arb_share_counter_next_value;
  wire             timer_1ms_s1_arb_share_set_values;
  wire             timer_1ms_s1_beginbursttransfer_internal;
  wire             timer_1ms_s1_begins_xfer;
  wire             timer_1ms_s1_chipselect;
  wire             timer_1ms_s1_end_xfer;
  wire             timer_1ms_s1_firsttransfer;
  wire             timer_1ms_s1_grant_vector;
  wire             timer_1ms_s1_in_a_read_cycle;
  wire             timer_1ms_s1_in_a_write_cycle;
  wire             timer_1ms_s1_irq_from_sa;
  wire             timer_1ms_s1_master_qreq_vector;
  wire             timer_1ms_s1_non_bursting_master_requests;
  wire    [ 15: 0] timer_1ms_s1_readdata_from_sa;
  reg              timer_1ms_s1_reg_firsttransfer;
  wire             timer_1ms_s1_reset_n;
  reg              timer_1ms_s1_slavearbiterlockenable;
  wire             timer_1ms_s1_slavearbiterlockenable2;
  wire             timer_1ms_s1_unreg_firsttransfer;
  wire             timer_1ms_s1_waits_for_read;
  wire             timer_1ms_s1_waits_for_write;
  wire             timer_1ms_s1_write_n;
  wire    [ 15: 0] timer_1ms_s1_writedata;
  wire             wait_for_timer_1ms_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~timer_1ms_s1_end_xfer;
    end


  assign timer_1ms_s1_begins_xfer = ~d1_reasons_to_wait & ((pb_cpu_to_io_m1_qualified_request_timer_1ms_s1));
  //assign timer_1ms_s1_readdata_from_sa = timer_1ms_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign timer_1ms_s1_readdata_from_sa = timer_1ms_s1_readdata;

  assign pb_cpu_to_io_m1_requests_timer_1ms_s1 = ({pb_cpu_to_io_m1_address_to_slave[22 : 5] , 5'b0} == 23'h400000) & pb_cpu_to_io_m1_chipselect;
  //timer_1ms_s1_arb_share_counter set values, which is an e_mux
  assign timer_1ms_s1_arb_share_set_values = 1;

  //timer_1ms_s1_non_bursting_master_requests mux, which is an e_mux
  assign timer_1ms_s1_non_bursting_master_requests = pb_cpu_to_io_m1_requests_timer_1ms_s1;

  //timer_1ms_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign timer_1ms_s1_any_bursting_master_saved_grant = 0;

  //timer_1ms_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign timer_1ms_s1_arb_share_counter_next_value = timer_1ms_s1_firsttransfer ? (timer_1ms_s1_arb_share_set_values - 1) : |timer_1ms_s1_arb_share_counter ? (timer_1ms_s1_arb_share_counter - 1) : 0;

  //timer_1ms_s1_allgrants all slave grants, which is an e_mux
  assign timer_1ms_s1_allgrants = |timer_1ms_s1_grant_vector;

  //timer_1ms_s1_end_xfer assignment, which is an e_assign
  assign timer_1ms_s1_end_xfer = ~(timer_1ms_s1_waits_for_read | timer_1ms_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_timer_1ms_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_timer_1ms_s1 = timer_1ms_s1_end_xfer & (~timer_1ms_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //timer_1ms_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign timer_1ms_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_timer_1ms_s1 & timer_1ms_s1_allgrants) | (end_xfer_arb_share_counter_term_timer_1ms_s1 & ~timer_1ms_s1_non_bursting_master_requests);

  //timer_1ms_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          timer_1ms_s1_arb_share_counter <= 0;
      else if (timer_1ms_s1_arb_counter_enable)
          timer_1ms_s1_arb_share_counter <= timer_1ms_s1_arb_share_counter_next_value;
    end


  //timer_1ms_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          timer_1ms_s1_slavearbiterlockenable <= 0;
      else if ((|timer_1ms_s1_master_qreq_vector & end_xfer_arb_share_counter_term_timer_1ms_s1) | (end_xfer_arb_share_counter_term_timer_1ms_s1 & ~timer_1ms_s1_non_bursting_master_requests))
          timer_1ms_s1_slavearbiterlockenable <= |timer_1ms_s1_arb_share_counter_next_value;
    end


  //pb_cpu_to_io/m1 timer_1ms/s1 arbiterlock, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock = timer_1ms_s1_slavearbiterlockenable & pb_cpu_to_io_m1_continuerequest;

  //timer_1ms_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign timer_1ms_s1_slavearbiterlockenable2 = |timer_1ms_s1_arb_share_counter_next_value;

  //pb_cpu_to_io/m1 timer_1ms/s1 arbiterlock2, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock2 = timer_1ms_s1_slavearbiterlockenable2 & pb_cpu_to_io_m1_continuerequest;

  //timer_1ms_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign timer_1ms_s1_any_continuerequest = 1;

  //pb_cpu_to_io_m1_continuerequest continued request, which is an e_assign
  assign pb_cpu_to_io_m1_continuerequest = 1;

  assign pb_cpu_to_io_m1_qualified_request_timer_1ms_s1 = pb_cpu_to_io_m1_requests_timer_1ms_s1 & ~(((pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ((pb_cpu_to_io_m1_latency_counter != 0))));
  //local readdatavalid pb_cpu_to_io_m1_read_data_valid_timer_1ms_s1, which is an e_mux
  assign pb_cpu_to_io_m1_read_data_valid_timer_1ms_s1 = pb_cpu_to_io_m1_granted_timer_1ms_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ~timer_1ms_s1_waits_for_read;

  //timer_1ms_s1_writedata mux, which is an e_mux
  assign timer_1ms_s1_writedata = pb_cpu_to_io_m1_writedata;

  //master is always granted when requested
  assign pb_cpu_to_io_m1_granted_timer_1ms_s1 = pb_cpu_to_io_m1_qualified_request_timer_1ms_s1;

  //pb_cpu_to_io/m1 saved-grant timer_1ms/s1, which is an e_assign
  assign pb_cpu_to_io_m1_saved_grant_timer_1ms_s1 = pb_cpu_to_io_m1_requests_timer_1ms_s1;

  //allow new arb cycle for timer_1ms/s1, which is an e_assign
  assign timer_1ms_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign timer_1ms_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign timer_1ms_s1_master_qreq_vector = 1;

  //timer_1ms_s1_reset_n assignment, which is an e_assign
  assign timer_1ms_s1_reset_n = reset_n;

  assign timer_1ms_s1_chipselect = pb_cpu_to_io_m1_granted_timer_1ms_s1;
  //timer_1ms_s1_firsttransfer first transaction, which is an e_assign
  assign timer_1ms_s1_firsttransfer = timer_1ms_s1_begins_xfer ? timer_1ms_s1_unreg_firsttransfer : timer_1ms_s1_reg_firsttransfer;

  //timer_1ms_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign timer_1ms_s1_unreg_firsttransfer = ~(timer_1ms_s1_slavearbiterlockenable & timer_1ms_s1_any_continuerequest);

  //timer_1ms_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          timer_1ms_s1_reg_firsttransfer <= 1'b1;
      else if (timer_1ms_s1_begins_xfer)
          timer_1ms_s1_reg_firsttransfer <= timer_1ms_s1_unreg_firsttransfer;
    end


  //timer_1ms_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign timer_1ms_s1_beginbursttransfer_internal = timer_1ms_s1_begins_xfer;

  //~timer_1ms_s1_write_n assignment, which is an e_mux
  assign timer_1ms_s1_write_n = ~(pb_cpu_to_io_m1_granted_timer_1ms_s1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect));

  assign shifted_address_to_timer_1ms_s1_from_pb_cpu_to_io_m1 = pb_cpu_to_io_m1_address_to_slave;
  //timer_1ms_s1_address mux, which is an e_mux
  assign timer_1ms_s1_address = shifted_address_to_timer_1ms_s1_from_pb_cpu_to_io_m1 >> 2;

  //d1_timer_1ms_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_timer_1ms_s1_end_xfer <= 1;
      else 
        d1_timer_1ms_s1_end_xfer <= timer_1ms_s1_end_xfer;
    end


  //timer_1ms_s1_waits_for_read in a cycle, which is an e_mux
  assign timer_1ms_s1_waits_for_read = timer_1ms_s1_in_a_read_cycle & timer_1ms_s1_begins_xfer;

  //timer_1ms_s1_in_a_read_cycle assignment, which is an e_assign
  assign timer_1ms_s1_in_a_read_cycle = pb_cpu_to_io_m1_granted_timer_1ms_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = timer_1ms_s1_in_a_read_cycle;

  //timer_1ms_s1_waits_for_write in a cycle, which is an e_mux
  assign timer_1ms_s1_waits_for_write = timer_1ms_s1_in_a_write_cycle & 0;

  //timer_1ms_s1_in_a_write_cycle assignment, which is an e_assign
  assign timer_1ms_s1_in_a_write_cycle = pb_cpu_to_io_m1_granted_timer_1ms_s1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = timer_1ms_s1_in_a_write_cycle;

  assign wait_for_timer_1ms_s1_counter = 0;
  //assign timer_1ms_s1_irq_from_sa = timer_1ms_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign timer_1ms_s1_irq_from_sa = timer_1ms_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //timer_1ms/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pb_cpu_to_io/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_io_m1_requests_timer_1ms_s1 && (pb_cpu_to_io_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pb_cpu_to_io/m1 drove 0 on its 'burstcount' port while accessing slave timer_1ms/s1", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tlb_miss_ram_1k_s1_arbitrator (
                                       // inputs:
                                        clk,
                                        cpu_tightly_coupled_instruction_master_0_address_to_slave,
                                        cpu_tightly_coupled_instruction_master_0_clken,
                                        cpu_tightly_coupled_instruction_master_0_latency_counter,
                                        cpu_tightly_coupled_instruction_master_0_read,
                                        reset_n,
                                        tlb_miss_ram_1k_s1_readdata,

                                       // outputs:
                                        cpu_tightly_coupled_instruction_master_0_granted_tlb_miss_ram_1k_s1,
                                        cpu_tightly_coupled_instruction_master_0_qualified_request_tlb_miss_ram_1k_s1,
                                        cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1,
                                        cpu_tightly_coupled_instruction_master_0_requests_tlb_miss_ram_1k_s1,
                                        d1_tlb_miss_ram_1k_s1_end_xfer,
                                        tlb_miss_ram_1k_s1_address,
                                        tlb_miss_ram_1k_s1_byteenable,
                                        tlb_miss_ram_1k_s1_chipselect,
                                        tlb_miss_ram_1k_s1_clken,
                                        tlb_miss_ram_1k_s1_readdata_from_sa,
                                        tlb_miss_ram_1k_s1_reset,
                                        tlb_miss_ram_1k_s1_write,
                                        tlb_miss_ram_1k_s1_writedata
                                     )
;

  output           cpu_tightly_coupled_instruction_master_0_granted_tlb_miss_ram_1k_s1;
  output           cpu_tightly_coupled_instruction_master_0_qualified_request_tlb_miss_ram_1k_s1;
  output           cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1;
  output           cpu_tightly_coupled_instruction_master_0_requests_tlb_miss_ram_1k_s1;
  output           d1_tlb_miss_ram_1k_s1_end_xfer;
  output  [  7: 0] tlb_miss_ram_1k_s1_address;
  output  [  3: 0] tlb_miss_ram_1k_s1_byteenable;
  output           tlb_miss_ram_1k_s1_chipselect;
  output           tlb_miss_ram_1k_s1_clken;
  output  [ 31: 0] tlb_miss_ram_1k_s1_readdata_from_sa;
  output           tlb_miss_ram_1k_s1_reset;
  output           tlb_miss_ram_1k_s1_write;
  output  [ 31: 0] tlb_miss_ram_1k_s1_writedata;
  input            clk;
  input   [ 26: 0] cpu_tightly_coupled_instruction_master_0_address_to_slave;
  input            cpu_tightly_coupled_instruction_master_0_clken;
  input            cpu_tightly_coupled_instruction_master_0_latency_counter;
  input            cpu_tightly_coupled_instruction_master_0_read;
  input            reset_n;
  input   [ 31: 0] tlb_miss_ram_1k_s1_readdata;

  wire             cpu_tightly_coupled_instruction_master_0_arbiterlock;
  wire             cpu_tightly_coupled_instruction_master_0_arbiterlock2;
  wire             cpu_tightly_coupled_instruction_master_0_continuerequest;
  wire             cpu_tightly_coupled_instruction_master_0_granted_tlb_miss_ram_1k_s1;
  wire             cpu_tightly_coupled_instruction_master_0_qualified_request_tlb_miss_ram_1k_s1;
  wire             cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1;
  reg              cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1_shift_register;
  wire             cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1_shift_register_in;
  wire             cpu_tightly_coupled_instruction_master_0_requests_tlb_miss_ram_1k_s1;
  wire             cpu_tightly_coupled_instruction_master_0_saved_grant_tlb_miss_ram_1k_s1;
  reg              d1_reasons_to_wait;
  reg              d1_tlb_miss_ram_1k_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_tlb_miss_ram_1k_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p1_cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1_shift_register;
  wire    [ 26: 0] shifted_address_to_tlb_miss_ram_1k_s1_from_cpu_tightly_coupled_instruction_master_0;
  wire    [  7: 0] tlb_miss_ram_1k_s1_address;
  wire             tlb_miss_ram_1k_s1_allgrants;
  wire             tlb_miss_ram_1k_s1_allow_new_arb_cycle;
  wire             tlb_miss_ram_1k_s1_any_bursting_master_saved_grant;
  wire             tlb_miss_ram_1k_s1_any_continuerequest;
  wire             tlb_miss_ram_1k_s1_arb_counter_enable;
  reg              tlb_miss_ram_1k_s1_arb_share_counter;
  wire             tlb_miss_ram_1k_s1_arb_share_counter_next_value;
  wire             tlb_miss_ram_1k_s1_arb_share_set_values;
  wire             tlb_miss_ram_1k_s1_beginbursttransfer_internal;
  wire             tlb_miss_ram_1k_s1_begins_xfer;
  wire    [  3: 0] tlb_miss_ram_1k_s1_byteenable;
  wire             tlb_miss_ram_1k_s1_chipselect;
  wire             tlb_miss_ram_1k_s1_clken;
  wire             tlb_miss_ram_1k_s1_end_xfer;
  wire             tlb_miss_ram_1k_s1_firsttransfer;
  wire             tlb_miss_ram_1k_s1_grant_vector;
  wire             tlb_miss_ram_1k_s1_in_a_read_cycle;
  wire             tlb_miss_ram_1k_s1_in_a_write_cycle;
  wire             tlb_miss_ram_1k_s1_master_qreq_vector;
  wire             tlb_miss_ram_1k_s1_non_bursting_master_requests;
  wire    [ 31: 0] tlb_miss_ram_1k_s1_readdata_from_sa;
  reg              tlb_miss_ram_1k_s1_reg_firsttransfer;
  wire             tlb_miss_ram_1k_s1_reset;
  reg              tlb_miss_ram_1k_s1_slavearbiterlockenable;
  wire             tlb_miss_ram_1k_s1_slavearbiterlockenable2;
  wire             tlb_miss_ram_1k_s1_unreg_firsttransfer;
  wire             tlb_miss_ram_1k_s1_waits_for_read;
  wire             tlb_miss_ram_1k_s1_waits_for_write;
  wire             tlb_miss_ram_1k_s1_write;
  wire    [ 31: 0] tlb_miss_ram_1k_s1_writedata;
  wire             wait_for_tlb_miss_ram_1k_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~tlb_miss_ram_1k_s1_end_xfer;
    end


  assign tlb_miss_ram_1k_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_tightly_coupled_instruction_master_0_qualified_request_tlb_miss_ram_1k_s1));
  //assign tlb_miss_ram_1k_s1_readdata_from_sa = tlb_miss_ram_1k_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tlb_miss_ram_1k_s1_readdata_from_sa = tlb_miss_ram_1k_s1_readdata;

  assign cpu_tightly_coupled_instruction_master_0_requests_tlb_miss_ram_1k_s1 = (({cpu_tightly_coupled_instruction_master_0_address_to_slave[26 : 10] , 10'b0} == 27'h7fff400) & (cpu_tightly_coupled_instruction_master_0_read)) & cpu_tightly_coupled_instruction_master_0_read;
  //tlb_miss_ram_1k_s1_arb_share_counter set values, which is an e_mux
  assign tlb_miss_ram_1k_s1_arb_share_set_values = 1;

  //tlb_miss_ram_1k_s1_non_bursting_master_requests mux, which is an e_mux
  assign tlb_miss_ram_1k_s1_non_bursting_master_requests = cpu_tightly_coupled_instruction_master_0_requests_tlb_miss_ram_1k_s1;

  //tlb_miss_ram_1k_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign tlb_miss_ram_1k_s1_any_bursting_master_saved_grant = 0;

  //tlb_miss_ram_1k_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign tlb_miss_ram_1k_s1_arb_share_counter_next_value = tlb_miss_ram_1k_s1_firsttransfer ? (tlb_miss_ram_1k_s1_arb_share_set_values - 1) : |tlb_miss_ram_1k_s1_arb_share_counter ? (tlb_miss_ram_1k_s1_arb_share_counter - 1) : 0;

  //tlb_miss_ram_1k_s1_allgrants all slave grants, which is an e_mux
  assign tlb_miss_ram_1k_s1_allgrants = |tlb_miss_ram_1k_s1_grant_vector;

  //tlb_miss_ram_1k_s1_end_xfer assignment, which is an e_assign
  assign tlb_miss_ram_1k_s1_end_xfer = ~(tlb_miss_ram_1k_s1_waits_for_read | tlb_miss_ram_1k_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_tlb_miss_ram_1k_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_tlb_miss_ram_1k_s1 = tlb_miss_ram_1k_s1_end_xfer & (~tlb_miss_ram_1k_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //tlb_miss_ram_1k_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign tlb_miss_ram_1k_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_tlb_miss_ram_1k_s1 & tlb_miss_ram_1k_s1_allgrants) | (end_xfer_arb_share_counter_term_tlb_miss_ram_1k_s1 & ~tlb_miss_ram_1k_s1_non_bursting_master_requests);

  //tlb_miss_ram_1k_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tlb_miss_ram_1k_s1_arb_share_counter <= 0;
      else if (tlb_miss_ram_1k_s1_arb_counter_enable)
          tlb_miss_ram_1k_s1_arb_share_counter <= tlb_miss_ram_1k_s1_arb_share_counter_next_value;
    end


  //tlb_miss_ram_1k_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tlb_miss_ram_1k_s1_slavearbiterlockenable <= 0;
      else if ((|tlb_miss_ram_1k_s1_master_qreq_vector & end_xfer_arb_share_counter_term_tlb_miss_ram_1k_s1) | (end_xfer_arb_share_counter_term_tlb_miss_ram_1k_s1 & ~tlb_miss_ram_1k_s1_non_bursting_master_requests))
          tlb_miss_ram_1k_s1_slavearbiterlockenable <= |tlb_miss_ram_1k_s1_arb_share_counter_next_value;
    end


  //cpu/tightly_coupled_instruction_master_0 tlb_miss_ram_1k/s1 arbiterlock, which is an e_assign
  assign cpu_tightly_coupled_instruction_master_0_arbiterlock = tlb_miss_ram_1k_s1_slavearbiterlockenable & cpu_tightly_coupled_instruction_master_0_continuerequest;

  //tlb_miss_ram_1k_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign tlb_miss_ram_1k_s1_slavearbiterlockenable2 = |tlb_miss_ram_1k_s1_arb_share_counter_next_value;

  //cpu/tightly_coupled_instruction_master_0 tlb_miss_ram_1k/s1 arbiterlock2, which is an e_assign
  assign cpu_tightly_coupled_instruction_master_0_arbiterlock2 = tlb_miss_ram_1k_s1_slavearbiterlockenable2 & cpu_tightly_coupled_instruction_master_0_continuerequest;

  //tlb_miss_ram_1k_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign tlb_miss_ram_1k_s1_any_continuerequest = 1;

  //cpu_tightly_coupled_instruction_master_0_continuerequest continued request, which is an e_assign
  assign cpu_tightly_coupled_instruction_master_0_continuerequest = 1;

  assign cpu_tightly_coupled_instruction_master_0_qualified_request_tlb_miss_ram_1k_s1 = cpu_tightly_coupled_instruction_master_0_requests_tlb_miss_ram_1k_s1;
  //cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1_shift_register_in = cpu_tightly_coupled_instruction_master_0_granted_tlb_miss_ram_1k_s1 & cpu_tightly_coupled_instruction_master_0_read & ~tlb_miss_ram_1k_s1_waits_for_read;

  //shift register p1 cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1_shift_register = {cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1_shift_register, cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1_shift_register_in};

  //cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1_shift_register <= 0;
      else 
        cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1_shift_register <= p1_cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1_shift_register;
    end


  //local readdatavalid cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1, which is an e_mux
  assign cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1 = cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1_shift_register;

  //mux tlb_miss_ram_1k_s1_clken, which is an e_mux
  assign tlb_miss_ram_1k_s1_clken = (cpu_tightly_coupled_instruction_master_0_granted_tlb_miss_ram_1k_s1)? cpu_tightly_coupled_instruction_master_0_clken :
    1'b1;

  //master is always granted when requested
  assign cpu_tightly_coupled_instruction_master_0_granted_tlb_miss_ram_1k_s1 = cpu_tightly_coupled_instruction_master_0_qualified_request_tlb_miss_ram_1k_s1;

  //cpu/tightly_coupled_instruction_master_0 saved-grant tlb_miss_ram_1k/s1, which is an e_assign
  assign cpu_tightly_coupled_instruction_master_0_saved_grant_tlb_miss_ram_1k_s1 = cpu_tightly_coupled_instruction_master_0_requests_tlb_miss_ram_1k_s1;

  //allow new arb cycle for tlb_miss_ram_1k/s1, which is an e_assign
  assign tlb_miss_ram_1k_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign tlb_miss_ram_1k_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign tlb_miss_ram_1k_s1_master_qreq_vector = 1;

  //~tlb_miss_ram_1k_s1_reset assignment, which is an e_assign
  assign tlb_miss_ram_1k_s1_reset = ~reset_n;

  assign tlb_miss_ram_1k_s1_chipselect = cpu_tightly_coupled_instruction_master_0_granted_tlb_miss_ram_1k_s1;
  //tlb_miss_ram_1k_s1_firsttransfer first transaction, which is an e_assign
  assign tlb_miss_ram_1k_s1_firsttransfer = tlb_miss_ram_1k_s1_begins_xfer ? tlb_miss_ram_1k_s1_unreg_firsttransfer : tlb_miss_ram_1k_s1_reg_firsttransfer;

  //tlb_miss_ram_1k_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign tlb_miss_ram_1k_s1_unreg_firsttransfer = ~(tlb_miss_ram_1k_s1_slavearbiterlockenable & tlb_miss_ram_1k_s1_any_continuerequest);

  //tlb_miss_ram_1k_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tlb_miss_ram_1k_s1_reg_firsttransfer <= 1'b1;
      else if (tlb_miss_ram_1k_s1_begins_xfer)
          tlb_miss_ram_1k_s1_reg_firsttransfer <= tlb_miss_ram_1k_s1_unreg_firsttransfer;
    end


  //tlb_miss_ram_1k_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign tlb_miss_ram_1k_s1_beginbursttransfer_internal = tlb_miss_ram_1k_s1_begins_xfer;

  //tlb_miss_ram_1k_s1_write assignment, which is an e_mux
  assign tlb_miss_ram_1k_s1_write = 0;

  assign shifted_address_to_tlb_miss_ram_1k_s1_from_cpu_tightly_coupled_instruction_master_0 = cpu_tightly_coupled_instruction_master_0_address_to_slave;
  //tlb_miss_ram_1k_s1_address mux, which is an e_mux
  assign tlb_miss_ram_1k_s1_address = shifted_address_to_tlb_miss_ram_1k_s1_from_cpu_tightly_coupled_instruction_master_0 >> 2;

  //d1_tlb_miss_ram_1k_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_tlb_miss_ram_1k_s1_end_xfer <= 1;
      else 
        d1_tlb_miss_ram_1k_s1_end_xfer <= tlb_miss_ram_1k_s1_end_xfer;
    end


  //tlb_miss_ram_1k_s1_waits_for_read in a cycle, which is an e_mux
  assign tlb_miss_ram_1k_s1_waits_for_read = tlb_miss_ram_1k_s1_in_a_read_cycle & 0;

  //tlb_miss_ram_1k_s1_in_a_read_cycle assignment, which is an e_assign
  assign tlb_miss_ram_1k_s1_in_a_read_cycle = cpu_tightly_coupled_instruction_master_0_granted_tlb_miss_ram_1k_s1 & cpu_tightly_coupled_instruction_master_0_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = tlb_miss_ram_1k_s1_in_a_read_cycle;

  //tlb_miss_ram_1k_s1_waits_for_write in a cycle, which is an e_mux
  assign tlb_miss_ram_1k_s1_waits_for_write = tlb_miss_ram_1k_s1_in_a_write_cycle & 0;

  //tlb_miss_ram_1k_s1_in_a_write_cycle assignment, which is an e_assign
  assign tlb_miss_ram_1k_s1_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = tlb_miss_ram_1k_s1_in_a_write_cycle;

  assign wait_for_tlb_miss_ram_1k_s1_counter = 0;
  //tlb_miss_ram_1k_s1_byteenable byte enable port mux, which is an e_mux
  assign tlb_miss_ram_1k_s1_byteenable = -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //tlb_miss_ram_1k/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tlb_miss_ram_1k_s2_arbitrator (
                                       // inputs:
                                        clk,
                                        cpu_tightly_coupled_data_master_0_address_to_slave,
                                        cpu_tightly_coupled_data_master_0_byteenable,
                                        cpu_tightly_coupled_data_master_0_clken,
                                        cpu_tightly_coupled_data_master_0_latency_counter,
                                        cpu_tightly_coupled_data_master_0_read,
                                        cpu_tightly_coupled_data_master_0_write,
                                        cpu_tightly_coupled_data_master_0_writedata,
                                        reset_n,
                                        tlb_miss_ram_1k_s2_readdata,

                                       // outputs:
                                        cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2,
                                        cpu_tightly_coupled_data_master_0_qualified_request_tlb_miss_ram_1k_s2,
                                        cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2,
                                        cpu_tightly_coupled_data_master_0_requests_tlb_miss_ram_1k_s2,
                                        d1_tlb_miss_ram_1k_s2_end_xfer,
                                        tlb_miss_ram_1k_s2_address,
                                        tlb_miss_ram_1k_s2_byteenable,
                                        tlb_miss_ram_1k_s2_chipselect,
                                        tlb_miss_ram_1k_s2_clken,
                                        tlb_miss_ram_1k_s2_readdata_from_sa,
                                        tlb_miss_ram_1k_s2_reset,
                                        tlb_miss_ram_1k_s2_write,
                                        tlb_miss_ram_1k_s2_writedata
                                     )
;

  output           cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2;
  output           cpu_tightly_coupled_data_master_0_qualified_request_tlb_miss_ram_1k_s2;
  output           cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2;
  output           cpu_tightly_coupled_data_master_0_requests_tlb_miss_ram_1k_s2;
  output           d1_tlb_miss_ram_1k_s2_end_xfer;
  output  [  7: 0] tlb_miss_ram_1k_s2_address;
  output  [  3: 0] tlb_miss_ram_1k_s2_byteenable;
  output           tlb_miss_ram_1k_s2_chipselect;
  output           tlb_miss_ram_1k_s2_clken;
  output  [ 31: 0] tlb_miss_ram_1k_s2_readdata_from_sa;
  output           tlb_miss_ram_1k_s2_reset;
  output           tlb_miss_ram_1k_s2_write;
  output  [ 31: 0] tlb_miss_ram_1k_s2_writedata;
  input            clk;
  input   [ 26: 0] cpu_tightly_coupled_data_master_0_address_to_slave;
  input   [  3: 0] cpu_tightly_coupled_data_master_0_byteenable;
  input            cpu_tightly_coupled_data_master_0_clken;
  input            cpu_tightly_coupled_data_master_0_latency_counter;
  input            cpu_tightly_coupled_data_master_0_read;
  input            cpu_tightly_coupled_data_master_0_write;
  input   [ 31: 0] cpu_tightly_coupled_data_master_0_writedata;
  input            reset_n;
  input   [ 31: 0] tlb_miss_ram_1k_s2_readdata;

  wire             cpu_tightly_coupled_data_master_0_arbiterlock;
  wire             cpu_tightly_coupled_data_master_0_arbiterlock2;
  wire             cpu_tightly_coupled_data_master_0_continuerequest;
  wire             cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2;
  wire             cpu_tightly_coupled_data_master_0_qualified_request_tlb_miss_ram_1k_s2;
  wire             cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2;
  reg              cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2_shift_register;
  wire             cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2_shift_register_in;
  wire             cpu_tightly_coupled_data_master_0_requests_tlb_miss_ram_1k_s2;
  wire             cpu_tightly_coupled_data_master_0_saved_grant_tlb_miss_ram_1k_s2;
  reg              d1_reasons_to_wait;
  reg              d1_tlb_miss_ram_1k_s2_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_tlb_miss_ram_1k_s2;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p1_cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2_shift_register;
  wire    [ 26: 0] shifted_address_to_tlb_miss_ram_1k_s2_from_cpu_tightly_coupled_data_master_0;
  wire    [  7: 0] tlb_miss_ram_1k_s2_address;
  wire             tlb_miss_ram_1k_s2_allgrants;
  wire             tlb_miss_ram_1k_s2_allow_new_arb_cycle;
  wire             tlb_miss_ram_1k_s2_any_bursting_master_saved_grant;
  wire             tlb_miss_ram_1k_s2_any_continuerequest;
  wire             tlb_miss_ram_1k_s2_arb_counter_enable;
  reg              tlb_miss_ram_1k_s2_arb_share_counter;
  wire             tlb_miss_ram_1k_s2_arb_share_counter_next_value;
  wire             tlb_miss_ram_1k_s2_arb_share_set_values;
  wire             tlb_miss_ram_1k_s2_beginbursttransfer_internal;
  wire             tlb_miss_ram_1k_s2_begins_xfer;
  wire    [  3: 0] tlb_miss_ram_1k_s2_byteenable;
  wire             tlb_miss_ram_1k_s2_chipselect;
  wire             tlb_miss_ram_1k_s2_clken;
  wire             tlb_miss_ram_1k_s2_end_xfer;
  wire             tlb_miss_ram_1k_s2_firsttransfer;
  wire             tlb_miss_ram_1k_s2_grant_vector;
  wire             tlb_miss_ram_1k_s2_in_a_read_cycle;
  wire             tlb_miss_ram_1k_s2_in_a_write_cycle;
  wire             tlb_miss_ram_1k_s2_master_qreq_vector;
  wire             tlb_miss_ram_1k_s2_non_bursting_master_requests;
  wire    [ 31: 0] tlb_miss_ram_1k_s2_readdata_from_sa;
  reg              tlb_miss_ram_1k_s2_reg_firsttransfer;
  wire             tlb_miss_ram_1k_s2_reset;
  reg              tlb_miss_ram_1k_s2_slavearbiterlockenable;
  wire             tlb_miss_ram_1k_s2_slavearbiterlockenable2;
  wire             tlb_miss_ram_1k_s2_unreg_firsttransfer;
  wire             tlb_miss_ram_1k_s2_waits_for_read;
  wire             tlb_miss_ram_1k_s2_waits_for_write;
  wire             tlb_miss_ram_1k_s2_write;
  wire    [ 31: 0] tlb_miss_ram_1k_s2_writedata;
  wire             wait_for_tlb_miss_ram_1k_s2_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~tlb_miss_ram_1k_s2_end_xfer;
    end


  assign tlb_miss_ram_1k_s2_begins_xfer = ~d1_reasons_to_wait & ((cpu_tightly_coupled_data_master_0_qualified_request_tlb_miss_ram_1k_s2));
  //assign tlb_miss_ram_1k_s2_readdata_from_sa = tlb_miss_ram_1k_s2_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tlb_miss_ram_1k_s2_readdata_from_sa = tlb_miss_ram_1k_s2_readdata;

  assign cpu_tightly_coupled_data_master_0_requests_tlb_miss_ram_1k_s2 = ({cpu_tightly_coupled_data_master_0_address_to_slave[26 : 10] , 10'b0} == 27'h7fff400) & (cpu_tightly_coupled_data_master_0_read | cpu_tightly_coupled_data_master_0_write);
  //tlb_miss_ram_1k_s2_arb_share_counter set values, which is an e_mux
  assign tlb_miss_ram_1k_s2_arb_share_set_values = 1;

  //tlb_miss_ram_1k_s2_non_bursting_master_requests mux, which is an e_mux
  assign tlb_miss_ram_1k_s2_non_bursting_master_requests = cpu_tightly_coupled_data_master_0_requests_tlb_miss_ram_1k_s2;

  //tlb_miss_ram_1k_s2_any_bursting_master_saved_grant mux, which is an e_mux
  assign tlb_miss_ram_1k_s2_any_bursting_master_saved_grant = 0;

  //tlb_miss_ram_1k_s2_arb_share_counter_next_value assignment, which is an e_assign
  assign tlb_miss_ram_1k_s2_arb_share_counter_next_value = tlb_miss_ram_1k_s2_firsttransfer ? (tlb_miss_ram_1k_s2_arb_share_set_values - 1) : |tlb_miss_ram_1k_s2_arb_share_counter ? (tlb_miss_ram_1k_s2_arb_share_counter - 1) : 0;

  //tlb_miss_ram_1k_s2_allgrants all slave grants, which is an e_mux
  assign tlb_miss_ram_1k_s2_allgrants = |tlb_miss_ram_1k_s2_grant_vector;

  //tlb_miss_ram_1k_s2_end_xfer assignment, which is an e_assign
  assign tlb_miss_ram_1k_s2_end_xfer = ~(tlb_miss_ram_1k_s2_waits_for_read | tlb_miss_ram_1k_s2_waits_for_write);

  //end_xfer_arb_share_counter_term_tlb_miss_ram_1k_s2 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_tlb_miss_ram_1k_s2 = tlb_miss_ram_1k_s2_end_xfer & (~tlb_miss_ram_1k_s2_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //tlb_miss_ram_1k_s2_arb_share_counter arbitration counter enable, which is an e_assign
  assign tlb_miss_ram_1k_s2_arb_counter_enable = (end_xfer_arb_share_counter_term_tlb_miss_ram_1k_s2 & tlb_miss_ram_1k_s2_allgrants) | (end_xfer_arb_share_counter_term_tlb_miss_ram_1k_s2 & ~tlb_miss_ram_1k_s2_non_bursting_master_requests);

  //tlb_miss_ram_1k_s2_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tlb_miss_ram_1k_s2_arb_share_counter <= 0;
      else if (tlb_miss_ram_1k_s2_arb_counter_enable)
          tlb_miss_ram_1k_s2_arb_share_counter <= tlb_miss_ram_1k_s2_arb_share_counter_next_value;
    end


  //tlb_miss_ram_1k_s2_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tlb_miss_ram_1k_s2_slavearbiterlockenable <= 0;
      else if ((|tlb_miss_ram_1k_s2_master_qreq_vector & end_xfer_arb_share_counter_term_tlb_miss_ram_1k_s2) | (end_xfer_arb_share_counter_term_tlb_miss_ram_1k_s2 & ~tlb_miss_ram_1k_s2_non_bursting_master_requests))
          tlb_miss_ram_1k_s2_slavearbiterlockenable <= |tlb_miss_ram_1k_s2_arb_share_counter_next_value;
    end


  //cpu/tightly_coupled_data_master_0 tlb_miss_ram_1k/s2 arbiterlock, which is an e_assign
  assign cpu_tightly_coupled_data_master_0_arbiterlock = tlb_miss_ram_1k_s2_slavearbiterlockenable & cpu_tightly_coupled_data_master_0_continuerequest;

  //tlb_miss_ram_1k_s2_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign tlb_miss_ram_1k_s2_slavearbiterlockenable2 = |tlb_miss_ram_1k_s2_arb_share_counter_next_value;

  //cpu/tightly_coupled_data_master_0 tlb_miss_ram_1k/s2 arbiterlock2, which is an e_assign
  assign cpu_tightly_coupled_data_master_0_arbiterlock2 = tlb_miss_ram_1k_s2_slavearbiterlockenable2 & cpu_tightly_coupled_data_master_0_continuerequest;

  //tlb_miss_ram_1k_s2_any_continuerequest at least one master continues requesting, which is an e_assign
  assign tlb_miss_ram_1k_s2_any_continuerequest = 1;

  //cpu_tightly_coupled_data_master_0_continuerequest continued request, which is an e_assign
  assign cpu_tightly_coupled_data_master_0_continuerequest = 1;

  assign cpu_tightly_coupled_data_master_0_qualified_request_tlb_miss_ram_1k_s2 = cpu_tightly_coupled_data_master_0_requests_tlb_miss_ram_1k_s2;
  //cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2_shift_register_in = cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2 & cpu_tightly_coupled_data_master_0_read & ~tlb_miss_ram_1k_s2_waits_for_read;

  //shift register p1 cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2_shift_register = {cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2_shift_register, cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2_shift_register_in};

  //cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2_shift_register <= 0;
      else 
        cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2_shift_register <= p1_cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2_shift_register;
    end


  //local readdatavalid cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2, which is an e_mux
  assign cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2 = cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2_shift_register;

  //tlb_miss_ram_1k_s2_writedata mux, which is an e_mux
  assign tlb_miss_ram_1k_s2_writedata = cpu_tightly_coupled_data_master_0_writedata;

  //mux tlb_miss_ram_1k_s2_clken, which is an e_mux
  assign tlb_miss_ram_1k_s2_clken = (cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2)? cpu_tightly_coupled_data_master_0_clken :
    1'b1;

  //master is always granted when requested
  assign cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2 = cpu_tightly_coupled_data_master_0_qualified_request_tlb_miss_ram_1k_s2;

  //cpu/tightly_coupled_data_master_0 saved-grant tlb_miss_ram_1k/s2, which is an e_assign
  assign cpu_tightly_coupled_data_master_0_saved_grant_tlb_miss_ram_1k_s2 = cpu_tightly_coupled_data_master_0_requests_tlb_miss_ram_1k_s2;

  //allow new arb cycle for tlb_miss_ram_1k/s2, which is an e_assign
  assign tlb_miss_ram_1k_s2_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign tlb_miss_ram_1k_s2_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign tlb_miss_ram_1k_s2_master_qreq_vector = 1;

  //~tlb_miss_ram_1k_s2_reset assignment, which is an e_assign
  assign tlb_miss_ram_1k_s2_reset = ~reset_n;

  assign tlb_miss_ram_1k_s2_chipselect = cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2;
  //tlb_miss_ram_1k_s2_firsttransfer first transaction, which is an e_assign
  assign tlb_miss_ram_1k_s2_firsttransfer = tlb_miss_ram_1k_s2_begins_xfer ? tlb_miss_ram_1k_s2_unreg_firsttransfer : tlb_miss_ram_1k_s2_reg_firsttransfer;

  //tlb_miss_ram_1k_s2_unreg_firsttransfer first transaction, which is an e_assign
  assign tlb_miss_ram_1k_s2_unreg_firsttransfer = ~(tlb_miss_ram_1k_s2_slavearbiterlockenable & tlb_miss_ram_1k_s2_any_continuerequest);

  //tlb_miss_ram_1k_s2_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tlb_miss_ram_1k_s2_reg_firsttransfer <= 1'b1;
      else if (tlb_miss_ram_1k_s2_begins_xfer)
          tlb_miss_ram_1k_s2_reg_firsttransfer <= tlb_miss_ram_1k_s2_unreg_firsttransfer;
    end


  //tlb_miss_ram_1k_s2_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign tlb_miss_ram_1k_s2_beginbursttransfer_internal = tlb_miss_ram_1k_s2_begins_xfer;

  //tlb_miss_ram_1k_s2_write assignment, which is an e_mux
  assign tlb_miss_ram_1k_s2_write = cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2 & cpu_tightly_coupled_data_master_0_write;

  assign shifted_address_to_tlb_miss_ram_1k_s2_from_cpu_tightly_coupled_data_master_0 = cpu_tightly_coupled_data_master_0_address_to_slave;
  //tlb_miss_ram_1k_s2_address mux, which is an e_mux
  assign tlb_miss_ram_1k_s2_address = shifted_address_to_tlb_miss_ram_1k_s2_from_cpu_tightly_coupled_data_master_0 >> 2;

  //d1_tlb_miss_ram_1k_s2_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_tlb_miss_ram_1k_s2_end_xfer <= 1;
      else 
        d1_tlb_miss_ram_1k_s2_end_xfer <= tlb_miss_ram_1k_s2_end_xfer;
    end


  //tlb_miss_ram_1k_s2_waits_for_read in a cycle, which is an e_mux
  assign tlb_miss_ram_1k_s2_waits_for_read = tlb_miss_ram_1k_s2_in_a_read_cycle & 0;

  //tlb_miss_ram_1k_s2_in_a_read_cycle assignment, which is an e_assign
  assign tlb_miss_ram_1k_s2_in_a_read_cycle = cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2 & cpu_tightly_coupled_data_master_0_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = tlb_miss_ram_1k_s2_in_a_read_cycle;

  //tlb_miss_ram_1k_s2_waits_for_write in a cycle, which is an e_mux
  assign tlb_miss_ram_1k_s2_waits_for_write = tlb_miss_ram_1k_s2_in_a_write_cycle & 0;

  //tlb_miss_ram_1k_s2_in_a_write_cycle assignment, which is an e_assign
  assign tlb_miss_ram_1k_s2_in_a_write_cycle = cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2 & cpu_tightly_coupled_data_master_0_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = tlb_miss_ram_1k_s2_in_a_write_cycle;

  assign wait_for_tlb_miss_ram_1k_s2_counter = 0;
  //tlb_miss_ram_1k_s2_byteenable byte enable port mux, which is an e_mux
  assign tlb_miss_ram_1k_s2_byteenable = (cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2)? cpu_tightly_coupled_data_master_0_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //tlb_miss_ram_1k/s2 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tse_mac_control_port_arbitrator (
                                         // inputs:
                                          clk,
                                          pb_cpu_to_io_m1_address_to_slave,
                                          pb_cpu_to_io_m1_burstcount,
                                          pb_cpu_to_io_m1_chipselect,
                                          pb_cpu_to_io_m1_latency_counter,
                                          pb_cpu_to_io_m1_read,
                                          pb_cpu_to_io_m1_write,
                                          pb_cpu_to_io_m1_writedata,
                                          reset_n,
                                          tse_mac_control_port_readdata,
                                          tse_mac_control_port_waitrequest,

                                         // outputs:
                                          d1_tse_mac_control_port_end_xfer,
                                          pb_cpu_to_io_m1_granted_tse_mac_control_port,
                                          pb_cpu_to_io_m1_qualified_request_tse_mac_control_port,
                                          pb_cpu_to_io_m1_read_data_valid_tse_mac_control_port,
                                          pb_cpu_to_io_m1_requests_tse_mac_control_port,
                                          tse_mac_control_port_address,
                                          tse_mac_control_port_read,
                                          tse_mac_control_port_readdata_from_sa,
                                          tse_mac_control_port_reset,
                                          tse_mac_control_port_waitrequest_from_sa,
                                          tse_mac_control_port_write,
                                          tse_mac_control_port_writedata
                                       )
;

  output           d1_tse_mac_control_port_end_xfer;
  output           pb_cpu_to_io_m1_granted_tse_mac_control_port;
  output           pb_cpu_to_io_m1_qualified_request_tse_mac_control_port;
  output           pb_cpu_to_io_m1_read_data_valid_tse_mac_control_port;
  output           pb_cpu_to_io_m1_requests_tse_mac_control_port;
  output  [  7: 0] tse_mac_control_port_address;
  output           tse_mac_control_port_read;
  output  [ 31: 0] tse_mac_control_port_readdata_from_sa;
  output           tse_mac_control_port_reset;
  output           tse_mac_control_port_waitrequest_from_sa;
  output           tse_mac_control_port_write;
  output  [ 31: 0] tse_mac_control_port_writedata;
  input            clk;
  input   [ 22: 0] pb_cpu_to_io_m1_address_to_slave;
  input            pb_cpu_to_io_m1_burstcount;
  input            pb_cpu_to_io_m1_chipselect;
  input            pb_cpu_to_io_m1_latency_counter;
  input            pb_cpu_to_io_m1_read;
  input            pb_cpu_to_io_m1_write;
  input   [ 31: 0] pb_cpu_to_io_m1_writedata;
  input            reset_n;
  input   [ 31: 0] tse_mac_control_port_readdata;
  input            tse_mac_control_port_waitrequest;

  reg              d1_reasons_to_wait;
  reg              d1_tse_mac_control_port_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_tse_mac_control_port;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             pb_cpu_to_io_m1_arbiterlock;
  wire             pb_cpu_to_io_m1_arbiterlock2;
  wire             pb_cpu_to_io_m1_continuerequest;
  wire             pb_cpu_to_io_m1_granted_tse_mac_control_port;
  wire             pb_cpu_to_io_m1_qualified_request_tse_mac_control_port;
  wire             pb_cpu_to_io_m1_read_data_valid_tse_mac_control_port;
  wire             pb_cpu_to_io_m1_requests_tse_mac_control_port;
  wire             pb_cpu_to_io_m1_saved_grant_tse_mac_control_port;
  wire    [ 22: 0] shifted_address_to_tse_mac_control_port_from_pb_cpu_to_io_m1;
  wire    [  7: 0] tse_mac_control_port_address;
  wire             tse_mac_control_port_allgrants;
  wire             tse_mac_control_port_allow_new_arb_cycle;
  wire             tse_mac_control_port_any_bursting_master_saved_grant;
  wire             tse_mac_control_port_any_continuerequest;
  wire             tse_mac_control_port_arb_counter_enable;
  reg              tse_mac_control_port_arb_share_counter;
  wire             tse_mac_control_port_arb_share_counter_next_value;
  wire             tse_mac_control_port_arb_share_set_values;
  wire             tse_mac_control_port_beginbursttransfer_internal;
  wire             tse_mac_control_port_begins_xfer;
  wire             tse_mac_control_port_end_xfer;
  wire             tse_mac_control_port_firsttransfer;
  wire             tse_mac_control_port_grant_vector;
  wire             tse_mac_control_port_in_a_read_cycle;
  wire             tse_mac_control_port_in_a_write_cycle;
  wire             tse_mac_control_port_master_qreq_vector;
  wire             tse_mac_control_port_non_bursting_master_requests;
  wire             tse_mac_control_port_read;
  wire    [ 31: 0] tse_mac_control_port_readdata_from_sa;
  reg              tse_mac_control_port_reg_firsttransfer;
  wire             tse_mac_control_port_reset;
  reg              tse_mac_control_port_slavearbiterlockenable;
  wire             tse_mac_control_port_slavearbiterlockenable2;
  wire             tse_mac_control_port_unreg_firsttransfer;
  wire             tse_mac_control_port_waitrequest_from_sa;
  wire             tse_mac_control_port_waits_for_read;
  wire             tse_mac_control_port_waits_for_write;
  wire             tse_mac_control_port_write;
  wire    [ 31: 0] tse_mac_control_port_writedata;
  wire             wait_for_tse_mac_control_port_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~tse_mac_control_port_end_xfer;
    end


  assign tse_mac_control_port_begins_xfer = ~d1_reasons_to_wait & ((pb_cpu_to_io_m1_qualified_request_tse_mac_control_port));
  //assign tse_mac_control_port_readdata_from_sa = tse_mac_control_port_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tse_mac_control_port_readdata_from_sa = tse_mac_control_port_readdata;

  assign pb_cpu_to_io_m1_requests_tse_mac_control_port = ({pb_cpu_to_io_m1_address_to_slave[22 : 10] , 10'b0} == 23'h4000) & pb_cpu_to_io_m1_chipselect;
  //assign tse_mac_control_port_waitrequest_from_sa = tse_mac_control_port_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tse_mac_control_port_waitrequest_from_sa = tse_mac_control_port_waitrequest;

  //tse_mac_control_port_arb_share_counter set values, which is an e_mux
  assign tse_mac_control_port_arb_share_set_values = 1;

  //tse_mac_control_port_non_bursting_master_requests mux, which is an e_mux
  assign tse_mac_control_port_non_bursting_master_requests = pb_cpu_to_io_m1_requests_tse_mac_control_port;

  //tse_mac_control_port_any_bursting_master_saved_grant mux, which is an e_mux
  assign tse_mac_control_port_any_bursting_master_saved_grant = 0;

  //tse_mac_control_port_arb_share_counter_next_value assignment, which is an e_assign
  assign tse_mac_control_port_arb_share_counter_next_value = tse_mac_control_port_firsttransfer ? (tse_mac_control_port_arb_share_set_values - 1) : |tse_mac_control_port_arb_share_counter ? (tse_mac_control_port_arb_share_counter - 1) : 0;

  //tse_mac_control_port_allgrants all slave grants, which is an e_mux
  assign tse_mac_control_port_allgrants = |tse_mac_control_port_grant_vector;

  //tse_mac_control_port_end_xfer assignment, which is an e_assign
  assign tse_mac_control_port_end_xfer = ~(tse_mac_control_port_waits_for_read | tse_mac_control_port_waits_for_write);

  //end_xfer_arb_share_counter_term_tse_mac_control_port arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_tse_mac_control_port = tse_mac_control_port_end_xfer & (~tse_mac_control_port_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //tse_mac_control_port_arb_share_counter arbitration counter enable, which is an e_assign
  assign tse_mac_control_port_arb_counter_enable = (end_xfer_arb_share_counter_term_tse_mac_control_port & tse_mac_control_port_allgrants) | (end_xfer_arb_share_counter_term_tse_mac_control_port & ~tse_mac_control_port_non_bursting_master_requests);

  //tse_mac_control_port_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tse_mac_control_port_arb_share_counter <= 0;
      else if (tse_mac_control_port_arb_counter_enable)
          tse_mac_control_port_arb_share_counter <= tse_mac_control_port_arb_share_counter_next_value;
    end


  //tse_mac_control_port_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tse_mac_control_port_slavearbiterlockenable <= 0;
      else if ((|tse_mac_control_port_master_qreq_vector & end_xfer_arb_share_counter_term_tse_mac_control_port) | (end_xfer_arb_share_counter_term_tse_mac_control_port & ~tse_mac_control_port_non_bursting_master_requests))
          tse_mac_control_port_slavearbiterlockenable <= |tse_mac_control_port_arb_share_counter_next_value;
    end


  //pb_cpu_to_io/m1 tse_mac/control_port arbiterlock, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock = tse_mac_control_port_slavearbiterlockenable & pb_cpu_to_io_m1_continuerequest;

  //tse_mac_control_port_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign tse_mac_control_port_slavearbiterlockenable2 = |tse_mac_control_port_arb_share_counter_next_value;

  //pb_cpu_to_io/m1 tse_mac/control_port arbiterlock2, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock2 = tse_mac_control_port_slavearbiterlockenable2 & pb_cpu_to_io_m1_continuerequest;

  //tse_mac_control_port_any_continuerequest at least one master continues requesting, which is an e_assign
  assign tse_mac_control_port_any_continuerequest = 1;

  //pb_cpu_to_io_m1_continuerequest continued request, which is an e_assign
  assign pb_cpu_to_io_m1_continuerequest = 1;

  assign pb_cpu_to_io_m1_qualified_request_tse_mac_control_port = pb_cpu_to_io_m1_requests_tse_mac_control_port & ~(((pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ((pb_cpu_to_io_m1_latency_counter != 0))));
  //local readdatavalid pb_cpu_to_io_m1_read_data_valid_tse_mac_control_port, which is an e_mux
  assign pb_cpu_to_io_m1_read_data_valid_tse_mac_control_port = pb_cpu_to_io_m1_granted_tse_mac_control_port & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ~tse_mac_control_port_waits_for_read;

  //tse_mac_control_port_writedata mux, which is an e_mux
  assign tse_mac_control_port_writedata = pb_cpu_to_io_m1_writedata;

  //master is always granted when requested
  assign pb_cpu_to_io_m1_granted_tse_mac_control_port = pb_cpu_to_io_m1_qualified_request_tse_mac_control_port;

  //pb_cpu_to_io/m1 saved-grant tse_mac/control_port, which is an e_assign
  assign pb_cpu_to_io_m1_saved_grant_tse_mac_control_port = pb_cpu_to_io_m1_requests_tse_mac_control_port;

  //allow new arb cycle for tse_mac/control_port, which is an e_assign
  assign tse_mac_control_port_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign tse_mac_control_port_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign tse_mac_control_port_master_qreq_vector = 1;

  //~tse_mac_control_port_reset assignment, which is an e_assign
  assign tse_mac_control_port_reset = ~reset_n;

  //tse_mac_control_port_firsttransfer first transaction, which is an e_assign
  assign tse_mac_control_port_firsttransfer = tse_mac_control_port_begins_xfer ? tse_mac_control_port_unreg_firsttransfer : tse_mac_control_port_reg_firsttransfer;

  //tse_mac_control_port_unreg_firsttransfer first transaction, which is an e_assign
  assign tse_mac_control_port_unreg_firsttransfer = ~(tse_mac_control_port_slavearbiterlockenable & tse_mac_control_port_any_continuerequest);

  //tse_mac_control_port_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tse_mac_control_port_reg_firsttransfer <= 1'b1;
      else if (tse_mac_control_port_begins_xfer)
          tse_mac_control_port_reg_firsttransfer <= tse_mac_control_port_unreg_firsttransfer;
    end


  //tse_mac_control_port_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign tse_mac_control_port_beginbursttransfer_internal = tse_mac_control_port_begins_xfer;

  //tse_mac_control_port_read assignment, which is an e_mux
  assign tse_mac_control_port_read = pb_cpu_to_io_m1_granted_tse_mac_control_port & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect);

  //tse_mac_control_port_write assignment, which is an e_mux
  assign tse_mac_control_port_write = pb_cpu_to_io_m1_granted_tse_mac_control_port & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect);

  assign shifted_address_to_tse_mac_control_port_from_pb_cpu_to_io_m1 = pb_cpu_to_io_m1_address_to_slave;
  //tse_mac_control_port_address mux, which is an e_mux
  assign tse_mac_control_port_address = shifted_address_to_tse_mac_control_port_from_pb_cpu_to_io_m1 >> 2;

  //d1_tse_mac_control_port_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_tse_mac_control_port_end_xfer <= 1;
      else 
        d1_tse_mac_control_port_end_xfer <= tse_mac_control_port_end_xfer;
    end


  //tse_mac_control_port_waits_for_read in a cycle, which is an e_mux
  assign tse_mac_control_port_waits_for_read = tse_mac_control_port_in_a_read_cycle & tse_mac_control_port_waitrequest_from_sa;

  //tse_mac_control_port_in_a_read_cycle assignment, which is an e_assign
  assign tse_mac_control_port_in_a_read_cycle = pb_cpu_to_io_m1_granted_tse_mac_control_port & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = tse_mac_control_port_in_a_read_cycle;

  //tse_mac_control_port_waits_for_write in a cycle, which is an e_mux
  assign tse_mac_control_port_waits_for_write = tse_mac_control_port_in_a_write_cycle & tse_mac_control_port_waitrequest_from_sa;

  //tse_mac_control_port_in_a_write_cycle assignment, which is an e_assign
  assign tse_mac_control_port_in_a_write_cycle = pb_cpu_to_io_m1_granted_tse_mac_control_port & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = tse_mac_control_port_in_a_write_cycle;

  assign wait_for_tse_mac_control_port_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //tse_mac/control_port enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pb_cpu_to_io/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_io_m1_requests_tse_mac_control_port && (pb_cpu_to_io_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pb_cpu_to_io/m1 drove 0 on its 'burstcount' port while accessing slave tse_mac/control_port", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tse_mac_transmit_arbitrator (
                                     // inputs:
                                      clk,
                                      reset_n,
                                      sgdma_tx_out_data,
                                      sgdma_tx_out_empty,
                                      sgdma_tx_out_endofpacket,
                                      sgdma_tx_out_error,
                                      sgdma_tx_out_startofpacket,
                                      sgdma_tx_out_valid,
                                      tse_mac_transmit_ready,

                                     // outputs:
                                      tse_mac_transmit_data,
                                      tse_mac_transmit_empty,
                                      tse_mac_transmit_endofpacket,
                                      tse_mac_transmit_error,
                                      tse_mac_transmit_ready_from_sa,
                                      tse_mac_transmit_startofpacket,
                                      tse_mac_transmit_valid
                                   )
;

  output  [ 31: 0] tse_mac_transmit_data;
  output  [  1: 0] tse_mac_transmit_empty;
  output           tse_mac_transmit_endofpacket;
  output           tse_mac_transmit_error;
  output           tse_mac_transmit_ready_from_sa;
  output           tse_mac_transmit_startofpacket;
  output           tse_mac_transmit_valid;
  input            clk;
  input            reset_n;
  input   [ 31: 0] sgdma_tx_out_data;
  input   [  1: 0] sgdma_tx_out_empty;
  input            sgdma_tx_out_endofpacket;
  input            sgdma_tx_out_error;
  input            sgdma_tx_out_startofpacket;
  input            sgdma_tx_out_valid;
  input            tse_mac_transmit_ready;

  wire    [ 31: 0] tse_mac_transmit_data;
  wire    [  1: 0] tse_mac_transmit_empty;
  wire             tse_mac_transmit_endofpacket;
  wire             tse_mac_transmit_error;
  wire             tse_mac_transmit_ready_from_sa;
  wire             tse_mac_transmit_startofpacket;
  wire             tse_mac_transmit_valid;
  //mux tse_mac_transmit_data, which is an e_mux
  assign tse_mac_transmit_data = sgdma_tx_out_data;

  //mux tse_mac_transmit_endofpacket, which is an e_mux
  assign tse_mac_transmit_endofpacket = sgdma_tx_out_endofpacket;

  //mux tse_mac_transmit_error, which is an e_mux
  assign tse_mac_transmit_error = sgdma_tx_out_error;

  //mux tse_mac_transmit_empty, which is an e_mux
  assign tse_mac_transmit_empty = sgdma_tx_out_empty;

  //assign tse_mac_transmit_ready_from_sa = tse_mac_transmit_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tse_mac_transmit_ready_from_sa = tse_mac_transmit_ready;

  //mux tse_mac_transmit_startofpacket, which is an e_mux
  assign tse_mac_transmit_startofpacket = sgdma_tx_out_startofpacket;

  //mux tse_mac_transmit_valid, which is an e_mux
  assign tse_mac_transmit_valid = sgdma_tx_out_valid;


endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tse_mac_receive_arbitrator (
                                    // inputs:
                                     clk,
                                     reset_n,
                                     sgdma_rx_in_ready_from_sa,
                                     tse_mac_receive_data,
                                     tse_mac_receive_empty,
                                     tse_mac_receive_endofpacket,
                                     tse_mac_receive_error,
                                     tse_mac_receive_startofpacket,
                                     tse_mac_receive_valid,

                                    // outputs:
                                     tse_mac_receive_ready
                                  )
;

  output           tse_mac_receive_ready;
  input            clk;
  input            reset_n;
  input            sgdma_rx_in_ready_from_sa;
  input   [ 31: 0] tse_mac_receive_data;
  input   [  1: 0] tse_mac_receive_empty;
  input            tse_mac_receive_endofpacket;
  input   [  5: 0] tse_mac_receive_error;
  input            tse_mac_receive_startofpacket;
  input            tse_mac_receive_valid;

  wire             tse_mac_receive_ready;
  //mux tse_mac_receive_ready, which is an e_mux
  assign tse_mac_receive_ready = sgdma_rx_in_ready_from_sa;


endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module uart_s1_arbitrator (
                            // inputs:
                             clk,
                             pb_cpu_to_io_m1_address_to_slave,
                             pb_cpu_to_io_m1_burstcount,
                             pb_cpu_to_io_m1_chipselect,
                             pb_cpu_to_io_m1_latency_counter,
                             pb_cpu_to_io_m1_read,
                             pb_cpu_to_io_m1_write,
                             pb_cpu_to_io_m1_writedata,
                             reset_n,
                             uart_s1_dataavailable,
                             uart_s1_irq,
                             uart_s1_readdata,
                             uart_s1_readyfordata,

                            // outputs:
                             d1_uart_s1_end_xfer,
                             pb_cpu_to_io_m1_granted_uart_s1,
                             pb_cpu_to_io_m1_qualified_request_uart_s1,
                             pb_cpu_to_io_m1_read_data_valid_uart_s1,
                             pb_cpu_to_io_m1_requests_uart_s1,
                             uart_s1_address,
                             uart_s1_begintransfer,
                             uart_s1_chipselect,
                             uart_s1_dataavailable_from_sa,
                             uart_s1_irq_from_sa,
                             uart_s1_read_n,
                             uart_s1_readdata_from_sa,
                             uart_s1_readyfordata_from_sa,
                             uart_s1_reset_n,
                             uart_s1_write_n,
                             uart_s1_writedata
                          )
;

  output           d1_uart_s1_end_xfer;
  output           pb_cpu_to_io_m1_granted_uart_s1;
  output           pb_cpu_to_io_m1_qualified_request_uart_s1;
  output           pb_cpu_to_io_m1_read_data_valid_uart_s1;
  output           pb_cpu_to_io_m1_requests_uart_s1;
  output  [  2: 0] uart_s1_address;
  output           uart_s1_begintransfer;
  output           uart_s1_chipselect;
  output           uart_s1_dataavailable_from_sa;
  output           uart_s1_irq_from_sa;
  output           uart_s1_read_n;
  output  [ 15: 0] uart_s1_readdata_from_sa;
  output           uart_s1_readyfordata_from_sa;
  output           uart_s1_reset_n;
  output           uart_s1_write_n;
  output  [ 15: 0] uart_s1_writedata;
  input            clk;
  input   [ 22: 0] pb_cpu_to_io_m1_address_to_slave;
  input            pb_cpu_to_io_m1_burstcount;
  input            pb_cpu_to_io_m1_chipselect;
  input            pb_cpu_to_io_m1_latency_counter;
  input            pb_cpu_to_io_m1_read;
  input            pb_cpu_to_io_m1_write;
  input   [ 31: 0] pb_cpu_to_io_m1_writedata;
  input            reset_n;
  input            uart_s1_dataavailable;
  input            uart_s1_irq;
  input   [ 15: 0] uart_s1_readdata;
  input            uart_s1_readyfordata;

  reg              d1_reasons_to_wait;
  reg              d1_uart_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_uart_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             pb_cpu_to_io_m1_arbiterlock;
  wire             pb_cpu_to_io_m1_arbiterlock2;
  wire             pb_cpu_to_io_m1_continuerequest;
  wire             pb_cpu_to_io_m1_granted_uart_s1;
  wire             pb_cpu_to_io_m1_qualified_request_uart_s1;
  wire             pb_cpu_to_io_m1_read_data_valid_uart_s1;
  wire             pb_cpu_to_io_m1_requests_uart_s1;
  wire             pb_cpu_to_io_m1_saved_grant_uart_s1;
  wire    [ 22: 0] shifted_address_to_uart_s1_from_pb_cpu_to_io_m1;
  wire    [  2: 0] uart_s1_address;
  wire             uart_s1_allgrants;
  wire             uart_s1_allow_new_arb_cycle;
  wire             uart_s1_any_bursting_master_saved_grant;
  wire             uart_s1_any_continuerequest;
  wire             uart_s1_arb_counter_enable;
  reg              uart_s1_arb_share_counter;
  wire             uart_s1_arb_share_counter_next_value;
  wire             uart_s1_arb_share_set_values;
  wire             uart_s1_beginbursttransfer_internal;
  wire             uart_s1_begins_xfer;
  wire             uart_s1_begintransfer;
  wire             uart_s1_chipselect;
  wire             uart_s1_dataavailable_from_sa;
  wire             uart_s1_end_xfer;
  wire             uart_s1_firsttransfer;
  wire             uart_s1_grant_vector;
  wire             uart_s1_in_a_read_cycle;
  wire             uart_s1_in_a_write_cycle;
  wire             uart_s1_irq_from_sa;
  wire             uart_s1_master_qreq_vector;
  wire             uart_s1_non_bursting_master_requests;
  wire             uart_s1_read_n;
  wire    [ 15: 0] uart_s1_readdata_from_sa;
  wire             uart_s1_readyfordata_from_sa;
  reg              uart_s1_reg_firsttransfer;
  wire             uart_s1_reset_n;
  reg              uart_s1_slavearbiterlockenable;
  wire             uart_s1_slavearbiterlockenable2;
  wire             uart_s1_unreg_firsttransfer;
  wire             uart_s1_waits_for_read;
  wire             uart_s1_waits_for_write;
  wire             uart_s1_write_n;
  wire    [ 15: 0] uart_s1_writedata;
  wire             wait_for_uart_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~uart_s1_end_xfer;
    end


  assign uart_s1_begins_xfer = ~d1_reasons_to_wait & ((pb_cpu_to_io_m1_qualified_request_uart_s1));
  //assign uart_s1_readdata_from_sa = uart_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign uart_s1_readdata_from_sa = uart_s1_readdata;

  assign pb_cpu_to_io_m1_requests_uart_s1 = ({pb_cpu_to_io_m1_address_to_slave[22 : 5] , 5'b0} == 23'h4c80) & pb_cpu_to_io_m1_chipselect;
  //assign uart_s1_dataavailable_from_sa = uart_s1_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign uart_s1_dataavailable_from_sa = uart_s1_dataavailable;

  //assign uart_s1_readyfordata_from_sa = uart_s1_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign uart_s1_readyfordata_from_sa = uart_s1_readyfordata;

  //uart_s1_arb_share_counter set values, which is an e_mux
  assign uart_s1_arb_share_set_values = 1;

  //uart_s1_non_bursting_master_requests mux, which is an e_mux
  assign uart_s1_non_bursting_master_requests = pb_cpu_to_io_m1_requests_uart_s1;

  //uart_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign uart_s1_any_bursting_master_saved_grant = 0;

  //uart_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign uart_s1_arb_share_counter_next_value = uart_s1_firsttransfer ? (uart_s1_arb_share_set_values - 1) : |uart_s1_arb_share_counter ? (uart_s1_arb_share_counter - 1) : 0;

  //uart_s1_allgrants all slave grants, which is an e_mux
  assign uart_s1_allgrants = |uart_s1_grant_vector;

  //uart_s1_end_xfer assignment, which is an e_assign
  assign uart_s1_end_xfer = ~(uart_s1_waits_for_read | uart_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_uart_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_uart_s1 = uart_s1_end_xfer & (~uart_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //uart_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign uart_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_uart_s1 & uart_s1_allgrants) | (end_xfer_arb_share_counter_term_uart_s1 & ~uart_s1_non_bursting_master_requests);

  //uart_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          uart_s1_arb_share_counter <= 0;
      else if (uart_s1_arb_counter_enable)
          uart_s1_arb_share_counter <= uart_s1_arb_share_counter_next_value;
    end


  //uart_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          uart_s1_slavearbiterlockenable <= 0;
      else if ((|uart_s1_master_qreq_vector & end_xfer_arb_share_counter_term_uart_s1) | (end_xfer_arb_share_counter_term_uart_s1 & ~uart_s1_non_bursting_master_requests))
          uart_s1_slavearbiterlockenable <= |uart_s1_arb_share_counter_next_value;
    end


  //pb_cpu_to_io/m1 uart/s1 arbiterlock, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock = uart_s1_slavearbiterlockenable & pb_cpu_to_io_m1_continuerequest;

  //uart_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign uart_s1_slavearbiterlockenable2 = |uart_s1_arb_share_counter_next_value;

  //pb_cpu_to_io/m1 uart/s1 arbiterlock2, which is an e_assign
  assign pb_cpu_to_io_m1_arbiterlock2 = uart_s1_slavearbiterlockenable2 & pb_cpu_to_io_m1_continuerequest;

  //uart_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign uart_s1_any_continuerequest = 1;

  //pb_cpu_to_io_m1_continuerequest continued request, which is an e_assign
  assign pb_cpu_to_io_m1_continuerequest = 1;

  assign pb_cpu_to_io_m1_qualified_request_uart_s1 = pb_cpu_to_io_m1_requests_uart_s1 & ~(((pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ((pb_cpu_to_io_m1_latency_counter != 0))));
  //local readdatavalid pb_cpu_to_io_m1_read_data_valid_uart_s1, which is an e_mux
  assign pb_cpu_to_io_m1_read_data_valid_uart_s1 = pb_cpu_to_io_m1_granted_uart_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect) & ~uart_s1_waits_for_read;

  //uart_s1_writedata mux, which is an e_mux
  assign uart_s1_writedata = pb_cpu_to_io_m1_writedata;

  //master is always granted when requested
  assign pb_cpu_to_io_m1_granted_uart_s1 = pb_cpu_to_io_m1_qualified_request_uart_s1;

  //pb_cpu_to_io/m1 saved-grant uart/s1, which is an e_assign
  assign pb_cpu_to_io_m1_saved_grant_uart_s1 = pb_cpu_to_io_m1_requests_uart_s1;

  //allow new arb cycle for uart/s1, which is an e_assign
  assign uart_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign uart_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign uart_s1_master_qreq_vector = 1;

  assign uart_s1_begintransfer = uart_s1_begins_xfer;
  //uart_s1_reset_n assignment, which is an e_assign
  assign uart_s1_reset_n = reset_n;

  assign uart_s1_chipselect = pb_cpu_to_io_m1_granted_uart_s1;
  //uart_s1_firsttransfer first transaction, which is an e_assign
  assign uart_s1_firsttransfer = uart_s1_begins_xfer ? uart_s1_unreg_firsttransfer : uart_s1_reg_firsttransfer;

  //uart_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign uart_s1_unreg_firsttransfer = ~(uart_s1_slavearbiterlockenable & uart_s1_any_continuerequest);

  //uart_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          uart_s1_reg_firsttransfer <= 1'b1;
      else if (uart_s1_begins_xfer)
          uart_s1_reg_firsttransfer <= uart_s1_unreg_firsttransfer;
    end


  //uart_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign uart_s1_beginbursttransfer_internal = uart_s1_begins_xfer;

  //~uart_s1_read_n assignment, which is an e_mux
  assign uart_s1_read_n = ~(pb_cpu_to_io_m1_granted_uart_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect));

  //~uart_s1_write_n assignment, which is an e_mux
  assign uart_s1_write_n = ~(pb_cpu_to_io_m1_granted_uart_s1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect));

  assign shifted_address_to_uart_s1_from_pb_cpu_to_io_m1 = pb_cpu_to_io_m1_address_to_slave;
  //uart_s1_address mux, which is an e_mux
  assign uart_s1_address = shifted_address_to_uart_s1_from_pb_cpu_to_io_m1 >> 2;

  //d1_uart_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_uart_s1_end_xfer <= 1;
      else 
        d1_uart_s1_end_xfer <= uart_s1_end_xfer;
    end


  //uart_s1_waits_for_read in a cycle, which is an e_mux
  assign uart_s1_waits_for_read = uart_s1_in_a_read_cycle & uart_s1_begins_xfer;

  //uart_s1_in_a_read_cycle assignment, which is an e_assign
  assign uart_s1_in_a_read_cycle = pb_cpu_to_io_m1_granted_uart_s1 & (pb_cpu_to_io_m1_read & pb_cpu_to_io_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = uart_s1_in_a_read_cycle;

  //uart_s1_waits_for_write in a cycle, which is an e_mux
  assign uart_s1_waits_for_write = uart_s1_in_a_write_cycle & uart_s1_begins_xfer;

  //uart_s1_in_a_write_cycle assignment, which is an e_assign
  assign uart_s1_in_a_write_cycle = pb_cpu_to_io_m1_granted_uart_s1 & (pb_cpu_to_io_m1_write & pb_cpu_to_io_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = uart_s1_in_a_write_cycle;

  assign wait_for_uart_s1_counter = 0;
  //assign uart_s1_irq_from_sa = uart_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign uart_s1_irq_from_sa = uart_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //uart/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pb_cpu_to_io/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pb_cpu_to_io_m1_requests_uart_s1 && (pb_cpu_to_io_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pb_cpu_to_io/m1 drove 0 on its 'burstcount' port while accessing slave uart/s1", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ghrd_4sgx230_sopc_reset_ddr3_top_phy_clk_out_domain_synch_module (
                                                                          // inputs:
                                                                           clk,
                                                                           data_in,
                                                                           reset_n,

                                                                          // outputs:
                                                                           data_out
                                                                        )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ghrd_4sgx230_sopc (
                           // 1) global signals:
                            clkin_100,
                            ddr3_top_aux_full_rate_clk_out,
                            ddr3_top_aux_half_rate_clk_out,
                            ddr3_top_phy_clk_out,
                            reset_n,

                           // the_button_pio
                            in_port_to_the_button_pio,

                           // the_ddr3_top
                            aux_scan_clk_from_the_ddr3_top,
                            aux_scan_clk_reset_n_from_the_ddr3_top,
                            dll_reference_clk_from_the_ddr3_top,
                            dqs_delay_ctrl_export_from_the_ddr3_top,
                            global_reset_n_to_the_ddr3_top,
                            local_init_done_from_the_ddr3_top,
                            local_refresh_ack_from_the_ddr3_top,
                            local_wdata_req_from_the_ddr3_top,
                            mem_addr_from_the_ddr3_top,
                            mem_ba_from_the_ddr3_top,
                            mem_cas_n_from_the_ddr3_top,
                            mem_cke_from_the_ddr3_top,
                            mem_clk_n_to_and_from_the_ddr3_top,
                            mem_clk_to_and_from_the_ddr3_top,
                            mem_cs_n_from_the_ddr3_top,
                            mem_dm_from_the_ddr3_top,
                            mem_dq_to_and_from_the_ddr3_top,
                            mem_dqs_to_and_from_the_ddr3_top,
                            mem_dqsn_to_and_from_the_ddr3_top,
                            mem_odt_from_the_ddr3_top,
                            mem_ras_n_from_the_ddr3_top,
                            mem_reset_n_from_the_ddr3_top,
                            mem_we_n_from_the_ddr3_top,
                            oct_ctl_rs_value_to_the_ddr3_top,
                            oct_ctl_rt_value_to_the_ddr3_top,
                            reset_phy_clk_n_from_the_ddr3_top,

                           // the_dipsw_pio
                            in_port_to_the_dipsw_pio,

                           // the_led_pio
                            out_port_from_the_led_pio,

                           // the_tb_fsm_avalon_slave
                            select_n_to_the_ext_flash,
                            select_n_to_the_ext_flash_1,
                            tb_fsm_address,
                            tb_fsm_data,
                            tb_fsm_readn,
                            tb_fsm_writen,

                           // the_tse_mac
                            led_an_from_the_tse_mac,
                            led_char_err_from_the_tse_mac,
                            led_col_from_the_tse_mac,
                            led_crs_from_the_tse_mac,
                            led_disp_err_from_the_tse_mac,
                            led_link_from_the_tse_mac,
                            mdc_from_the_tse_mac,
                            mdio_in_to_the_tse_mac,
                            mdio_oen_from_the_tse_mac,
                            mdio_out_from_the_tse_mac,
                            ref_clk_to_the_tse_mac,
                            rx_recovclkout_from_the_tse_mac,
                            rxp_to_the_tse_mac,
                            txp_from_the_tse_mac,

                           // the_uart
                            rxd_to_the_uart,
                            txd_from_the_uart
                         )
;

  output           aux_scan_clk_from_the_ddr3_top;
  output           aux_scan_clk_reset_n_from_the_ddr3_top;
  output           ddr3_top_aux_full_rate_clk_out;
  output           ddr3_top_aux_half_rate_clk_out;
  output           ddr3_top_phy_clk_out;
  output           dll_reference_clk_from_the_ddr3_top;
  output  [  5: 0] dqs_delay_ctrl_export_from_the_ddr3_top;
  output           led_an_from_the_tse_mac;
  output           led_char_err_from_the_tse_mac;
  output           led_col_from_the_tse_mac;
  output           led_crs_from_the_tse_mac;
  output           led_disp_err_from_the_tse_mac;
  output           led_link_from_the_tse_mac;
  output           local_init_done_from_the_ddr3_top;
  output           local_refresh_ack_from_the_ddr3_top;
  output           local_wdata_req_from_the_ddr3_top;
  output           mdc_from_the_tse_mac;
  output           mdio_oen_from_the_tse_mac;
  output           mdio_out_from_the_tse_mac;
  output  [ 12: 0] mem_addr_from_the_ddr3_top;
  output  [  2: 0] mem_ba_from_the_ddr3_top;
  output           mem_cas_n_from_the_ddr3_top;
  output           mem_cke_from_the_ddr3_top;
  inout            mem_clk_n_to_and_from_the_ddr3_top;
  inout            mem_clk_to_and_from_the_ddr3_top;
  output           mem_cs_n_from_the_ddr3_top;
  output  [  1: 0] mem_dm_from_the_ddr3_top;
  inout   [ 15: 0] mem_dq_to_and_from_the_ddr3_top;
  inout   [  1: 0] mem_dqs_to_and_from_the_ddr3_top;
  inout   [  1: 0] mem_dqsn_to_and_from_the_ddr3_top;
  output           mem_odt_from_the_ddr3_top;
  output           mem_ras_n_from_the_ddr3_top;
  output           mem_reset_n_from_the_ddr3_top;
  output           mem_we_n_from_the_ddr3_top;
  output  [ 15: 0] out_port_from_the_led_pio;
  output           reset_phy_clk_n_from_the_ddr3_top;
  output           rx_recovclkout_from_the_tse_mac;
  output           select_n_to_the_ext_flash;
  output           select_n_to_the_ext_flash_1;
  output  [ 24: 0] tb_fsm_address;
  inout   [ 15: 0] tb_fsm_data;
  output           tb_fsm_readn;
  output           tb_fsm_writen;
  output           txd_from_the_uart;
  output           txp_from_the_tse_mac;
  input            clkin_100;
  input            global_reset_n_to_the_ddr3_top;
  input   [  2: 0] in_port_to_the_button_pio;
  input   [  7: 0] in_port_to_the_dipsw_pio;
  input            mdio_in_to_the_tse_mac;
  input   [ 13: 0] oct_ctl_rs_value_to_the_ddr3_top;
  input   [ 13: 0] oct_ctl_rt_value_to_the_ddr3_top;
  input            ref_clk_to_the_tse_mac;
  input            reset_n;
  input            rxd_to_the_uart;
  input            rxp_to_the_tse_mac;

  wire             aux_scan_clk_from_the_ddr3_top;
  wire             aux_scan_clk_reset_n_from_the_ddr3_top;
  wire    [  1: 0] button_pio_s1_address;
  wire             button_pio_s1_chipselect;
  wire             button_pio_s1_irq;
  wire             button_pio_s1_irq_from_sa;
  wire    [  2: 0] button_pio_s1_readdata;
  wire    [  2: 0] button_pio_s1_readdata_from_sa;
  wire             button_pio_s1_reset_n;
  wire             button_pio_s1_write_n;
  wire    [  2: 0] button_pio_s1_writedata;
  wire             clkin_100_reset_n;
  wire    [ 28: 0] cpu_data_master_address;
  wire    [ 28: 0] cpu_data_master_address_to_slave;
  wire    [  3: 0] cpu_data_master_byteenable;
  wire             cpu_data_master_debugaccess;
  wire             cpu_data_master_granted_cpu_jtag_debug_module;
  wire             cpu_data_master_granted_pb_cpu_to_ddr3_top_s1;
  wire             cpu_data_master_granted_pb_cpu_to_fsm_s1;
  wire             cpu_data_master_granted_pb_cpu_to_io_s1;
  wire    [ 31: 0] cpu_data_master_irq;
  wire             cpu_data_master_latency_counter;
  wire             cpu_data_master_qualified_request_cpu_jtag_debug_module;
  wire             cpu_data_master_qualified_request_pb_cpu_to_ddr3_top_s1;
  wire             cpu_data_master_qualified_request_pb_cpu_to_fsm_s1;
  wire             cpu_data_master_qualified_request_pb_cpu_to_io_s1;
  wire             cpu_data_master_read;
  wire             cpu_data_master_read_data_valid_cpu_jtag_debug_module;
  wire             cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1;
  wire             cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register;
  wire             cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1;
  wire             cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register;
  wire             cpu_data_master_read_data_valid_pb_cpu_to_io_s1;
  wire             cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register;
  wire    [ 31: 0] cpu_data_master_readdata;
  wire             cpu_data_master_readdatavalid;
  wire             cpu_data_master_requests_cpu_jtag_debug_module;
  wire             cpu_data_master_requests_pb_cpu_to_ddr3_top_s1;
  wire             cpu_data_master_requests_pb_cpu_to_fsm_s1;
  wire             cpu_data_master_requests_pb_cpu_to_io_s1;
  wire             cpu_data_master_waitrequest;
  wire             cpu_data_master_write;
  wire    [ 31: 0] cpu_data_master_writedata;
  wire    [ 28: 0] cpu_instruction_master_address;
  wire    [ 28: 0] cpu_instruction_master_address_to_slave;
  wire             cpu_instruction_master_granted_cpu_jtag_debug_module;
  wire             cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1;
  wire             cpu_instruction_master_granted_pb_cpu_to_fsm_s1;
  wire             cpu_instruction_master_latency_counter;
  wire             cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  wire             cpu_instruction_master_qualified_request_pb_cpu_to_ddr3_top_s1;
  wire             cpu_instruction_master_qualified_request_pb_cpu_to_fsm_s1;
  wire             cpu_instruction_master_read;
  wire             cpu_instruction_master_read_data_valid_cpu_jtag_debug_module;
  wire             cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1;
  wire             cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register;
  wire             cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1;
  wire             cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register;
  wire    [ 31: 0] cpu_instruction_master_readdata;
  wire             cpu_instruction_master_readdatavalid;
  wire             cpu_instruction_master_requests_cpu_jtag_debug_module;
  wire             cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1;
  wire             cpu_instruction_master_requests_pb_cpu_to_fsm_s1;
  wire             cpu_instruction_master_waitrequest;
  wire    [  8: 0] cpu_jtag_debug_module_address;
  wire             cpu_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_jtag_debug_module_byteenable;
  wire             cpu_jtag_debug_module_chipselect;
  wire             cpu_jtag_debug_module_debugaccess;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  wire             cpu_jtag_debug_module_reset_n;
  wire             cpu_jtag_debug_module_resetrequest;
  wire             cpu_jtag_debug_module_resetrequest_from_sa;
  wire             cpu_jtag_debug_module_write;
  wire    [ 31: 0] cpu_jtag_debug_module_writedata;
  wire    [ 26: 0] cpu_tightly_coupled_data_master_0_address;
  wire    [ 26: 0] cpu_tightly_coupled_data_master_0_address_to_slave;
  wire    [  3: 0] cpu_tightly_coupled_data_master_0_byteenable;
  wire             cpu_tightly_coupled_data_master_0_clken;
  wire             cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2;
  wire             cpu_tightly_coupled_data_master_0_latency_counter;
  wire             cpu_tightly_coupled_data_master_0_qualified_request_tlb_miss_ram_1k_s2;
  wire             cpu_tightly_coupled_data_master_0_read;
  wire             cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2;
  wire    [ 31: 0] cpu_tightly_coupled_data_master_0_readdata;
  wire             cpu_tightly_coupled_data_master_0_readdatavalid;
  wire             cpu_tightly_coupled_data_master_0_requests_tlb_miss_ram_1k_s2;
  wire             cpu_tightly_coupled_data_master_0_waitrequest;
  wire             cpu_tightly_coupled_data_master_0_write;
  wire    [ 31: 0] cpu_tightly_coupled_data_master_0_writedata;
  wire    [ 26: 0] cpu_tightly_coupled_instruction_master_0_address;
  wire    [ 26: 0] cpu_tightly_coupled_instruction_master_0_address_to_slave;
  wire             cpu_tightly_coupled_instruction_master_0_clken;
  wire             cpu_tightly_coupled_instruction_master_0_granted_tlb_miss_ram_1k_s1;
  wire             cpu_tightly_coupled_instruction_master_0_latency_counter;
  wire             cpu_tightly_coupled_instruction_master_0_qualified_request_tlb_miss_ram_1k_s1;
  wire             cpu_tightly_coupled_instruction_master_0_read;
  wire             cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1;
  wire    [ 31: 0] cpu_tightly_coupled_instruction_master_0_readdata;
  wire             cpu_tightly_coupled_instruction_master_0_readdatavalid;
  wire             cpu_tightly_coupled_instruction_master_0_requests_tlb_miss_ram_1k_s1;
  wire             cpu_tightly_coupled_instruction_master_0_waitrequest;
  wire             d1_button_pio_s1_end_xfer;
  wire             d1_cpu_jtag_debug_module_end_xfer;
  wire             d1_ddr3_top_s1_end_xfer;
  wire             d1_descriptor_memory_s1_end_xfer;
  wire             d1_dipsw_pio_s1_end_xfer;
  wire             d1_jtag_uart_avalon_jtag_slave_end_xfer;
  wire             d1_led_pio_s1_end_xfer;
  wire             d1_pb_cpu_to_ddr3_top_s1_end_xfer;
  wire             d1_pb_cpu_to_fsm_s1_end_xfer;
  wire             d1_pb_cpu_to_io_s1_end_xfer;
  wire             d1_pb_dma_to_ddr3_top_s1_end_xfer;
  wire             d1_pb_dma_to_descriptor_memory_s1_end_xfer;
  wire             d1_sgdma_rx_csr_end_xfer;
  wire             d1_sgdma_tx_csr_end_xfer;
  wire             d1_sysid_control_slave_end_xfer;
  wire             d1_tb_fsm_avalon_slave_end_xfer;
  wire             d1_timer_1ms_s1_end_xfer;
  wire             d1_tlb_miss_ram_1k_s1_end_xfer;
  wire             d1_tlb_miss_ram_1k_s2_end_xfer;
  wire             d1_tse_mac_control_port_end_xfer;
  wire             d1_uart_s1_end_xfer;
  wire             ddr3_top_aux_full_rate_clk_out;
  wire             ddr3_top_aux_half_rate_clk_out;
  wire             ddr3_top_phy_clk_out;
  wire             ddr3_top_phy_clk_out_reset_n;
  wire    [ 23: 0] ddr3_top_s1_address;
  wire             ddr3_top_s1_beginbursttransfer;
  wire    [  2: 0] ddr3_top_s1_burstcount;
  wire    [  7: 0] ddr3_top_s1_byteenable;
  wire             ddr3_top_s1_read;
  wire    [ 63: 0] ddr3_top_s1_readdata;
  wire    [ 63: 0] ddr3_top_s1_readdata_from_sa;
  wire             ddr3_top_s1_readdatavalid;
  wire             ddr3_top_s1_resetrequest_n;
  wire             ddr3_top_s1_resetrequest_n_from_sa;
  wire             ddr3_top_s1_waitrequest_n;
  wire             ddr3_top_s1_waitrequest_n_from_sa;
  wire             ddr3_top_s1_write;
  wire    [ 63: 0] ddr3_top_s1_writedata;
  wire    [ 10: 0] descriptor_memory_s1_address;
  wire    [  3: 0] descriptor_memory_s1_byteenable;
  wire             descriptor_memory_s1_chipselect;
  wire             descriptor_memory_s1_clken;
  wire    [ 31: 0] descriptor_memory_s1_readdata;
  wire    [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  wire             descriptor_memory_s1_reset;
  wire             descriptor_memory_s1_write;
  wire    [ 31: 0] descriptor_memory_s1_writedata;
  wire    [  1: 0] dipsw_pio_s1_address;
  wire             dipsw_pio_s1_chipselect;
  wire             dipsw_pio_s1_irq;
  wire             dipsw_pio_s1_irq_from_sa;
  wire    [  7: 0] dipsw_pio_s1_readdata;
  wire    [  7: 0] dipsw_pio_s1_readdata_from_sa;
  wire             dipsw_pio_s1_reset_n;
  wire             dipsw_pio_s1_write_n;
  wire    [  7: 0] dipsw_pio_s1_writedata;
  wire             dll_reference_clk_from_the_ddr3_top;
  wire    [  5: 0] dqs_delay_ctrl_export_from_the_ddr3_top;
  wire             ext_flash_1_s1_wait_counter_eq_0;
  wire             ext_flash_s1_wait_counter_eq_0;
  wire    [ 15: 0] incoming_tb_fsm_data_with_Xs_converted_to_0;
  wire             jtag_uart_avalon_jtag_slave_address;
  wire             jtag_uart_avalon_jtag_slave_chipselect;
  wire             jtag_uart_avalon_jtag_slave_dataavailable;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_irq;
  wire             jtag_uart_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_reset_n;
  wire             jtag_uart_avalon_jtag_slave_waitrequest;
  wire             jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  wire             led_an_from_the_tse_mac;
  wire             led_char_err_from_the_tse_mac;
  wire             led_col_from_the_tse_mac;
  wire             led_crs_from_the_tse_mac;
  wire             led_disp_err_from_the_tse_mac;
  wire             led_link_from_the_tse_mac;
  wire    [  1: 0] led_pio_s1_address;
  wire             led_pio_s1_chipselect;
  wire    [ 15: 0] led_pio_s1_readdata;
  wire    [ 15: 0] led_pio_s1_readdata_from_sa;
  wire             led_pio_s1_reset_n;
  wire             led_pio_s1_write_n;
  wire    [ 15: 0] led_pio_s1_writedata;
  wire             local_init_done_from_the_ddr3_top;
  wire             local_refresh_ack_from_the_ddr3_top;
  wire             local_wdata_req_from_the_ddr3_top;
  wire             mdc_from_the_tse_mac;
  wire             mdio_oen_from_the_tse_mac;
  wire             mdio_out_from_the_tse_mac;
  wire    [ 12: 0] mem_addr_from_the_ddr3_top;
  wire    [  2: 0] mem_ba_from_the_ddr3_top;
  wire             mem_cas_n_from_the_ddr3_top;
  wire             mem_cke_from_the_ddr3_top;
  wire             mem_clk_n_to_and_from_the_ddr3_top;
  wire             mem_clk_to_and_from_the_ddr3_top;
  wire             mem_cs_n_from_the_ddr3_top;
  wire    [  1: 0] mem_dm_from_the_ddr3_top;
  wire    [ 15: 0] mem_dq_to_and_from_the_ddr3_top;
  wire    [  1: 0] mem_dqs_to_and_from_the_ddr3_top;
  wire    [  1: 0] mem_dqsn_to_and_from_the_ddr3_top;
  wire             mem_odt_from_the_ddr3_top;
  wire             mem_ras_n_from_the_ddr3_top;
  wire             mem_reset_n_from_the_ddr3_top;
  wire             mem_we_n_from_the_ddr3_top;
  wire             out_clk_ddr3_top_aux_full_rate_clk;
  wire             out_clk_ddr3_top_aux_half_rate_clk;
  wire             out_clk_ddr3_top_phy_clk;
  wire    [ 15: 0] out_port_from_the_led_pio;
  wire    [ 26: 0] pb_cpu_to_ddr3_top_m1_address;
  wire    [ 26: 0] pb_cpu_to_ddr3_top_m1_address_to_slave;
  wire             pb_cpu_to_ddr3_top_m1_burstcount;
  wire    [  3: 0] pb_cpu_to_ddr3_top_m1_byteenable;
  wire             pb_cpu_to_ddr3_top_m1_chipselect;
  wire             pb_cpu_to_ddr3_top_m1_debugaccess;
  wire             pb_cpu_to_ddr3_top_m1_endofpacket;
  wire             pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1;
  wire             pb_cpu_to_ddr3_top_m1_latency_counter;
  wire             pb_cpu_to_ddr3_top_m1_qualified_request_ddr3_top_s1;
  wire             pb_cpu_to_ddr3_top_m1_read;
  wire             pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1;
  wire             pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register;
  wire    [ 31: 0] pb_cpu_to_ddr3_top_m1_readdata;
  wire             pb_cpu_to_ddr3_top_m1_readdatavalid;
  wire             pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1;
  wire             pb_cpu_to_ddr3_top_m1_waitrequest;
  wire             pb_cpu_to_ddr3_top_m1_write;
  wire    [ 31: 0] pb_cpu_to_ddr3_top_m1_writedata;
  wire    [ 24: 0] pb_cpu_to_ddr3_top_s1_address;
  wire             pb_cpu_to_ddr3_top_s1_arbiterlock;
  wire             pb_cpu_to_ddr3_top_s1_arbiterlock2;
  wire             pb_cpu_to_ddr3_top_s1_burstcount;
  wire    [  3: 0] pb_cpu_to_ddr3_top_s1_byteenable;
  wire             pb_cpu_to_ddr3_top_s1_chipselect;
  wire             pb_cpu_to_ddr3_top_s1_debugaccess;
  wire             pb_cpu_to_ddr3_top_s1_endofpacket;
  wire             pb_cpu_to_ddr3_top_s1_endofpacket_from_sa;
  wire    [ 24: 0] pb_cpu_to_ddr3_top_s1_nativeaddress;
  wire             pb_cpu_to_ddr3_top_s1_read;
  wire    [ 31: 0] pb_cpu_to_ddr3_top_s1_readdata;
  wire    [ 31: 0] pb_cpu_to_ddr3_top_s1_readdata_from_sa;
  wire             pb_cpu_to_ddr3_top_s1_readdatavalid;
  wire             pb_cpu_to_ddr3_top_s1_reset_n;
  wire             pb_cpu_to_ddr3_top_s1_waitrequest;
  wire             pb_cpu_to_ddr3_top_s1_waitrequest_from_sa;
  wire             pb_cpu_to_ddr3_top_s1_write;
  wire    [ 31: 0] pb_cpu_to_ddr3_top_s1_writedata;
  wire    [ 25: 0] pb_cpu_to_fsm_m1_address;
  wire    [ 25: 0] pb_cpu_to_fsm_m1_address_to_slave;
  wire             pb_cpu_to_fsm_m1_burstcount;
  wire    [  3: 0] pb_cpu_to_fsm_m1_byteenable;
  wire    [  1: 0] pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1;
  wire    [  1: 0] pb_cpu_to_fsm_m1_byteenable_ext_flash_s1;
  wire             pb_cpu_to_fsm_m1_chipselect;
  wire    [  1: 0] pb_cpu_to_fsm_m1_dbs_address;
  wire    [ 15: 0] pb_cpu_to_fsm_m1_dbs_write_16;
  wire             pb_cpu_to_fsm_m1_debugaccess;
  wire             pb_cpu_to_fsm_m1_endofpacket;
  wire             pb_cpu_to_fsm_m1_granted_ext_flash_1_s1;
  wire             pb_cpu_to_fsm_m1_granted_ext_flash_s1;
  wire    [  1: 0] pb_cpu_to_fsm_m1_latency_counter;
  wire             pb_cpu_to_fsm_m1_qualified_request_ext_flash_1_s1;
  wire             pb_cpu_to_fsm_m1_qualified_request_ext_flash_s1;
  wire             pb_cpu_to_fsm_m1_read;
  wire             pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1;
  wire             pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1;
  wire    [ 31: 0] pb_cpu_to_fsm_m1_readdata;
  wire             pb_cpu_to_fsm_m1_readdatavalid;
  wire             pb_cpu_to_fsm_m1_requests_ext_flash_1_s1;
  wire             pb_cpu_to_fsm_m1_requests_ext_flash_s1;
  wire             pb_cpu_to_fsm_m1_waitrequest;
  wire             pb_cpu_to_fsm_m1_write;
  wire    [ 31: 0] pb_cpu_to_fsm_m1_writedata;
  wire    [ 23: 0] pb_cpu_to_fsm_s1_address;
  wire             pb_cpu_to_fsm_s1_arbiterlock;
  wire             pb_cpu_to_fsm_s1_arbiterlock2;
  wire             pb_cpu_to_fsm_s1_burstcount;
  wire    [  3: 0] pb_cpu_to_fsm_s1_byteenable;
  wire             pb_cpu_to_fsm_s1_chipselect;
  wire             pb_cpu_to_fsm_s1_debugaccess;
  wire             pb_cpu_to_fsm_s1_endofpacket;
  wire             pb_cpu_to_fsm_s1_endofpacket_from_sa;
  wire    [ 23: 0] pb_cpu_to_fsm_s1_nativeaddress;
  wire             pb_cpu_to_fsm_s1_read;
  wire    [ 31: 0] pb_cpu_to_fsm_s1_readdata;
  wire    [ 31: 0] pb_cpu_to_fsm_s1_readdata_from_sa;
  wire             pb_cpu_to_fsm_s1_readdatavalid;
  wire             pb_cpu_to_fsm_s1_reset_n;
  wire             pb_cpu_to_fsm_s1_waitrequest;
  wire             pb_cpu_to_fsm_s1_waitrequest_from_sa;
  wire             pb_cpu_to_fsm_s1_write;
  wire    [ 31: 0] pb_cpu_to_fsm_s1_writedata;
  wire    [ 22: 0] pb_cpu_to_io_m1_address;
  wire    [ 22: 0] pb_cpu_to_io_m1_address_to_slave;
  wire             pb_cpu_to_io_m1_burstcount;
  wire    [  3: 0] pb_cpu_to_io_m1_byteenable;
  wire             pb_cpu_to_io_m1_chipselect;
  wire             pb_cpu_to_io_m1_debugaccess;
  wire             pb_cpu_to_io_m1_endofpacket;
  wire             pb_cpu_to_io_m1_granted_button_pio_s1;
  wire             pb_cpu_to_io_m1_granted_descriptor_memory_s1;
  wire             pb_cpu_to_io_m1_granted_dipsw_pio_s1;
  wire             pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave;
  wire             pb_cpu_to_io_m1_granted_led_pio_s1;
  wire             pb_cpu_to_io_m1_granted_sgdma_rx_csr;
  wire             pb_cpu_to_io_m1_granted_sgdma_tx_csr;
  wire             pb_cpu_to_io_m1_granted_sysid_control_slave;
  wire             pb_cpu_to_io_m1_granted_timer_1ms_s1;
  wire             pb_cpu_to_io_m1_granted_tse_mac_control_port;
  wire             pb_cpu_to_io_m1_granted_uart_s1;
  wire             pb_cpu_to_io_m1_latency_counter;
  wire             pb_cpu_to_io_m1_qualified_request_button_pio_s1;
  wire             pb_cpu_to_io_m1_qualified_request_descriptor_memory_s1;
  wire             pb_cpu_to_io_m1_qualified_request_dipsw_pio_s1;
  wire             pb_cpu_to_io_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  wire             pb_cpu_to_io_m1_qualified_request_led_pio_s1;
  wire             pb_cpu_to_io_m1_qualified_request_sgdma_rx_csr;
  wire             pb_cpu_to_io_m1_qualified_request_sgdma_tx_csr;
  wire             pb_cpu_to_io_m1_qualified_request_sysid_control_slave;
  wire             pb_cpu_to_io_m1_qualified_request_timer_1ms_s1;
  wire             pb_cpu_to_io_m1_qualified_request_tse_mac_control_port;
  wire             pb_cpu_to_io_m1_qualified_request_uart_s1;
  wire             pb_cpu_to_io_m1_read;
  wire             pb_cpu_to_io_m1_read_data_valid_button_pio_s1;
  wire             pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1;
  wire             pb_cpu_to_io_m1_read_data_valid_dipsw_pio_s1;
  wire             pb_cpu_to_io_m1_read_data_valid_jtag_uart_avalon_jtag_slave;
  wire             pb_cpu_to_io_m1_read_data_valid_led_pio_s1;
  wire             pb_cpu_to_io_m1_read_data_valid_sgdma_rx_csr;
  wire             pb_cpu_to_io_m1_read_data_valid_sgdma_tx_csr;
  wire             pb_cpu_to_io_m1_read_data_valid_sysid_control_slave;
  wire             pb_cpu_to_io_m1_read_data_valid_timer_1ms_s1;
  wire             pb_cpu_to_io_m1_read_data_valid_tse_mac_control_port;
  wire             pb_cpu_to_io_m1_read_data_valid_uart_s1;
  wire    [ 31: 0] pb_cpu_to_io_m1_readdata;
  wire             pb_cpu_to_io_m1_readdatavalid;
  wire             pb_cpu_to_io_m1_requests_button_pio_s1;
  wire             pb_cpu_to_io_m1_requests_descriptor_memory_s1;
  wire             pb_cpu_to_io_m1_requests_dipsw_pio_s1;
  wire             pb_cpu_to_io_m1_requests_jtag_uart_avalon_jtag_slave;
  wire             pb_cpu_to_io_m1_requests_led_pio_s1;
  wire             pb_cpu_to_io_m1_requests_sgdma_rx_csr;
  wire             pb_cpu_to_io_m1_requests_sgdma_tx_csr;
  wire             pb_cpu_to_io_m1_requests_sysid_control_slave;
  wire             pb_cpu_to_io_m1_requests_timer_1ms_s1;
  wire             pb_cpu_to_io_m1_requests_tse_mac_control_port;
  wire             pb_cpu_to_io_m1_requests_uart_s1;
  wire             pb_cpu_to_io_m1_waitrequest;
  wire             pb_cpu_to_io_m1_write;
  wire    [ 31: 0] pb_cpu_to_io_m1_writedata;
  wire    [ 20: 0] pb_cpu_to_io_s1_address;
  wire             pb_cpu_to_io_s1_arbiterlock;
  wire             pb_cpu_to_io_s1_arbiterlock2;
  wire             pb_cpu_to_io_s1_burstcount;
  wire    [  3: 0] pb_cpu_to_io_s1_byteenable;
  wire             pb_cpu_to_io_s1_chipselect;
  wire             pb_cpu_to_io_s1_debugaccess;
  wire             pb_cpu_to_io_s1_endofpacket;
  wire             pb_cpu_to_io_s1_endofpacket_from_sa;
  wire    [ 20: 0] pb_cpu_to_io_s1_nativeaddress;
  wire             pb_cpu_to_io_s1_read;
  wire    [ 31: 0] pb_cpu_to_io_s1_readdata;
  wire    [ 31: 0] pb_cpu_to_io_s1_readdata_from_sa;
  wire             pb_cpu_to_io_s1_readdatavalid;
  wire             pb_cpu_to_io_s1_reset_n;
  wire             pb_cpu_to_io_s1_waitrequest;
  wire             pb_cpu_to_io_s1_waitrequest_from_sa;
  wire             pb_cpu_to_io_s1_write;
  wire    [ 31: 0] pb_cpu_to_io_s1_writedata;
  wire    [ 26: 0] pb_dma_to_ddr3_top_m1_address;
  wire    [ 26: 0] pb_dma_to_ddr3_top_m1_address_to_slave;
  wire             pb_dma_to_ddr3_top_m1_burstcount;
  wire    [  3: 0] pb_dma_to_ddr3_top_m1_byteenable;
  wire             pb_dma_to_ddr3_top_m1_chipselect;
  wire             pb_dma_to_ddr3_top_m1_debugaccess;
  wire             pb_dma_to_ddr3_top_m1_endofpacket;
  wire             pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1;
  wire             pb_dma_to_ddr3_top_m1_latency_counter;
  wire             pb_dma_to_ddr3_top_m1_qualified_request_ddr3_top_s1;
  wire             pb_dma_to_ddr3_top_m1_read;
  wire             pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1;
  wire             pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register;
  wire    [ 31: 0] pb_dma_to_ddr3_top_m1_readdata;
  wire             pb_dma_to_ddr3_top_m1_readdatavalid;
  wire             pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1;
  wire             pb_dma_to_ddr3_top_m1_waitrequest;
  wire             pb_dma_to_ddr3_top_m1_write;
  wire    [ 31: 0] pb_dma_to_ddr3_top_m1_writedata;
  wire    [ 24: 0] pb_dma_to_ddr3_top_s1_address;
  wire             pb_dma_to_ddr3_top_s1_arbiterlock;
  wire             pb_dma_to_ddr3_top_s1_arbiterlock2;
  wire             pb_dma_to_ddr3_top_s1_burstcount;
  wire    [  3: 0] pb_dma_to_ddr3_top_s1_byteenable;
  wire             pb_dma_to_ddr3_top_s1_chipselect;
  wire             pb_dma_to_ddr3_top_s1_debugaccess;
  wire             pb_dma_to_ddr3_top_s1_endofpacket;
  wire             pb_dma_to_ddr3_top_s1_endofpacket_from_sa;
  wire    [ 24: 0] pb_dma_to_ddr3_top_s1_nativeaddress;
  wire             pb_dma_to_ddr3_top_s1_read;
  wire    [ 31: 0] pb_dma_to_ddr3_top_s1_readdata;
  wire    [ 31: 0] pb_dma_to_ddr3_top_s1_readdata_from_sa;
  wire             pb_dma_to_ddr3_top_s1_readdatavalid;
  wire             pb_dma_to_ddr3_top_s1_reset_n;
  wire             pb_dma_to_ddr3_top_s1_waitrequest;
  wire             pb_dma_to_ddr3_top_s1_waitrequest_from_sa;
  wire             pb_dma_to_ddr3_top_s1_write;
  wire    [ 31: 0] pb_dma_to_ddr3_top_s1_writedata;
  wire    [ 13: 0] pb_dma_to_descriptor_memory_m1_address;
  wire    [ 13: 0] pb_dma_to_descriptor_memory_m1_address_to_slave;
  wire             pb_dma_to_descriptor_memory_m1_burstcount;
  wire    [  3: 0] pb_dma_to_descriptor_memory_m1_byteenable;
  wire             pb_dma_to_descriptor_memory_m1_chipselect;
  wire             pb_dma_to_descriptor_memory_m1_debugaccess;
  wire             pb_dma_to_descriptor_memory_m1_endofpacket;
  wire             pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1;
  wire             pb_dma_to_descriptor_memory_m1_latency_counter;
  wire             pb_dma_to_descriptor_memory_m1_qualified_request_descriptor_memory_s1;
  wire             pb_dma_to_descriptor_memory_m1_read;
  wire             pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1;
  wire    [ 31: 0] pb_dma_to_descriptor_memory_m1_readdata;
  wire             pb_dma_to_descriptor_memory_m1_readdatavalid;
  wire             pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1;
  wire             pb_dma_to_descriptor_memory_m1_waitrequest;
  wire             pb_dma_to_descriptor_memory_m1_write;
  wire    [ 31: 0] pb_dma_to_descriptor_memory_m1_writedata;
  wire    [ 11: 0] pb_dma_to_descriptor_memory_s1_address;
  wire             pb_dma_to_descriptor_memory_s1_arbiterlock;
  wire             pb_dma_to_descriptor_memory_s1_arbiterlock2;
  wire             pb_dma_to_descriptor_memory_s1_burstcount;
  wire    [  3: 0] pb_dma_to_descriptor_memory_s1_byteenable;
  wire             pb_dma_to_descriptor_memory_s1_chipselect;
  wire             pb_dma_to_descriptor_memory_s1_debugaccess;
  wire             pb_dma_to_descriptor_memory_s1_endofpacket;
  wire             pb_dma_to_descriptor_memory_s1_endofpacket_from_sa;
  wire    [ 11: 0] pb_dma_to_descriptor_memory_s1_nativeaddress;
  wire             pb_dma_to_descriptor_memory_s1_read;
  wire    [ 31: 0] pb_dma_to_descriptor_memory_s1_readdata;
  wire    [ 31: 0] pb_dma_to_descriptor_memory_s1_readdata_from_sa;
  wire             pb_dma_to_descriptor_memory_s1_readdatavalid;
  wire             pb_dma_to_descriptor_memory_s1_reset_n;
  wire             pb_dma_to_descriptor_memory_s1_waitrequest;
  wire             pb_dma_to_descriptor_memory_s1_waitrequest_from_sa;
  wire             pb_dma_to_descriptor_memory_s1_write;
  wire    [ 31: 0] pb_dma_to_descriptor_memory_s1_writedata;
  wire             reset_n_sources;
  wire             reset_phy_clk_n_from_the_ddr3_top;
  wire             rx_recovclkout_from_the_tse_mac;
  wire             select_n_to_the_ext_flash;
  wire             select_n_to_the_ext_flash_1;
  wire    [  3: 0] sgdma_rx_csr_address;
  wire             sgdma_rx_csr_chipselect;
  wire             sgdma_rx_csr_irq;
  wire             sgdma_rx_csr_irq_from_sa;
  wire             sgdma_rx_csr_read;
  wire    [ 31: 0] sgdma_rx_csr_readdata;
  wire    [ 31: 0] sgdma_rx_csr_readdata_from_sa;
  wire             sgdma_rx_csr_reset_n;
  wire             sgdma_rx_csr_write;
  wire    [ 31: 0] sgdma_rx_csr_writedata;
  wire    [ 31: 0] sgdma_rx_descriptor_read_address;
  wire    [ 31: 0] sgdma_rx_descriptor_read_address_to_slave;
  wire             sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_latency_counter;
  wire             sgdma_rx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_read;
  wire             sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register;
  wire    [ 31: 0] sgdma_rx_descriptor_read_readdata;
  wire             sgdma_rx_descriptor_read_readdatavalid;
  wire             sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_waitrequest;
  wire    [ 31: 0] sgdma_rx_descriptor_write_address;
  wire    [ 31: 0] sgdma_rx_descriptor_write_address_to_slave;
  wire             sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_waitrequest;
  wire             sgdma_rx_descriptor_write_write;
  wire    [ 31: 0] sgdma_rx_descriptor_write_writedata;
  wire    [ 31: 0] sgdma_rx_in_data;
  wire    [  1: 0] sgdma_rx_in_empty;
  wire             sgdma_rx_in_endofpacket;
  wire    [  5: 0] sgdma_rx_in_error;
  wire             sgdma_rx_in_ready;
  wire             sgdma_rx_in_ready_from_sa;
  wire             sgdma_rx_in_startofpacket;
  wire             sgdma_rx_in_valid;
  wire    [ 31: 0] sgdma_rx_m_write_address;
  wire    [ 31: 0] sgdma_rx_m_write_address_to_slave;
  wire    [  3: 0] sgdma_rx_m_write_byteenable;
  wire             sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1;
  wire             sgdma_rx_m_write_qualified_request_pb_dma_to_ddr3_top_s1;
  wire             sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1;
  wire             sgdma_rx_m_write_waitrequest;
  wire             sgdma_rx_m_write_write;
  wire    [ 31: 0] sgdma_rx_m_write_writedata;
  wire    [  3: 0] sgdma_tx_csr_address;
  wire             sgdma_tx_csr_chipselect;
  wire             sgdma_tx_csr_irq;
  wire             sgdma_tx_csr_irq_from_sa;
  wire             sgdma_tx_csr_read;
  wire    [ 31: 0] sgdma_tx_csr_readdata;
  wire    [ 31: 0] sgdma_tx_csr_readdata_from_sa;
  wire             sgdma_tx_csr_reset_n;
  wire             sgdma_tx_csr_write;
  wire    [ 31: 0] sgdma_tx_csr_writedata;
  wire    [ 31: 0] sgdma_tx_descriptor_read_address;
  wire    [ 31: 0] sgdma_tx_descriptor_read_address_to_slave;
  wire             sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_latency_counter;
  wire             sgdma_tx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_read;
  wire             sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register;
  wire    [ 31: 0] sgdma_tx_descriptor_read_readdata;
  wire             sgdma_tx_descriptor_read_readdatavalid;
  wire             sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_waitrequest;
  wire    [ 31: 0] sgdma_tx_descriptor_write_address;
  wire    [ 31: 0] sgdma_tx_descriptor_write_address_to_slave;
  wire             sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_waitrequest;
  wire             sgdma_tx_descriptor_write_write;
  wire    [ 31: 0] sgdma_tx_descriptor_write_writedata;
  wire    [ 31: 0] sgdma_tx_m_read_address;
  wire    [ 31: 0] sgdma_tx_m_read_address_to_slave;
  wire             sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1;
  wire             sgdma_tx_m_read_latency_counter;
  wire             sgdma_tx_m_read_qualified_request_pb_dma_to_ddr3_top_s1;
  wire             sgdma_tx_m_read_read;
  wire             sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1;
  wire             sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1_shift_register;
  wire    [ 31: 0] sgdma_tx_m_read_readdata;
  wire             sgdma_tx_m_read_readdatavalid;
  wire             sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1;
  wire             sgdma_tx_m_read_waitrequest;
  wire    [ 31: 0] sgdma_tx_out_data;
  wire    [  1: 0] sgdma_tx_out_empty;
  wire             sgdma_tx_out_endofpacket;
  wire             sgdma_tx_out_error;
  wire             sgdma_tx_out_ready;
  wire             sgdma_tx_out_startofpacket;
  wire             sgdma_tx_out_valid;
  wire             sysid_control_slave_address;
  wire             sysid_control_slave_clock;
  wire    [ 31: 0] sysid_control_slave_readdata;
  wire    [ 31: 0] sysid_control_slave_readdata_from_sa;
  wire             sysid_control_slave_reset_n;
  wire    [ 24: 0] tb_fsm_address;
  wire    [ 15: 0] tb_fsm_data;
  wire             tb_fsm_readn;
  wire             tb_fsm_writen;
  wire    [  2: 0] timer_1ms_s1_address;
  wire             timer_1ms_s1_chipselect;
  wire             timer_1ms_s1_irq;
  wire             timer_1ms_s1_irq_from_sa;
  wire    [ 15: 0] timer_1ms_s1_readdata;
  wire    [ 15: 0] timer_1ms_s1_readdata_from_sa;
  wire             timer_1ms_s1_reset_n;
  wire             timer_1ms_s1_write_n;
  wire    [ 15: 0] timer_1ms_s1_writedata;
  wire    [  7: 0] tlb_miss_ram_1k_s1_address;
  wire    [  3: 0] tlb_miss_ram_1k_s1_byteenable;
  wire             tlb_miss_ram_1k_s1_chipselect;
  wire             tlb_miss_ram_1k_s1_clken;
  wire    [ 31: 0] tlb_miss_ram_1k_s1_readdata;
  wire    [ 31: 0] tlb_miss_ram_1k_s1_readdata_from_sa;
  wire             tlb_miss_ram_1k_s1_reset;
  wire             tlb_miss_ram_1k_s1_write;
  wire    [ 31: 0] tlb_miss_ram_1k_s1_writedata;
  wire    [  7: 0] tlb_miss_ram_1k_s2_address;
  wire    [  3: 0] tlb_miss_ram_1k_s2_byteenable;
  wire             tlb_miss_ram_1k_s2_chipselect;
  wire             tlb_miss_ram_1k_s2_clken;
  wire    [ 31: 0] tlb_miss_ram_1k_s2_readdata;
  wire    [ 31: 0] tlb_miss_ram_1k_s2_readdata_from_sa;
  wire             tlb_miss_ram_1k_s2_reset;
  wire             tlb_miss_ram_1k_s2_write;
  wire    [ 31: 0] tlb_miss_ram_1k_s2_writedata;
  wire    [  7: 0] tse_mac_control_port_address;
  wire             tse_mac_control_port_read;
  wire    [ 31: 0] tse_mac_control_port_readdata;
  wire    [ 31: 0] tse_mac_control_port_readdata_from_sa;
  wire             tse_mac_control_port_reset;
  wire             tse_mac_control_port_waitrequest;
  wire             tse_mac_control_port_waitrequest_from_sa;
  wire             tse_mac_control_port_write;
  wire    [ 31: 0] tse_mac_control_port_writedata;
  wire    [ 31: 0] tse_mac_receive_data;
  wire    [  1: 0] tse_mac_receive_empty;
  wire             tse_mac_receive_endofpacket;
  wire    [  5: 0] tse_mac_receive_error;
  wire             tse_mac_receive_ready;
  wire             tse_mac_receive_startofpacket;
  wire             tse_mac_receive_valid;
  wire    [ 31: 0] tse_mac_transmit_data;
  wire    [  1: 0] tse_mac_transmit_empty;
  wire             tse_mac_transmit_endofpacket;
  wire             tse_mac_transmit_error;
  wire             tse_mac_transmit_ready;
  wire             tse_mac_transmit_ready_from_sa;
  wire             tse_mac_transmit_startofpacket;
  wire             tse_mac_transmit_valid;
  wire             txd_from_the_uart;
  wire             txp_from_the_tse_mac;
  wire    [  2: 0] uart_s1_address;
  wire             uart_s1_begintransfer;
  wire             uart_s1_chipselect;
  wire             uart_s1_dataavailable;
  wire             uart_s1_dataavailable_from_sa;
  wire             uart_s1_irq;
  wire             uart_s1_irq_from_sa;
  wire             uart_s1_read_n;
  wire    [ 15: 0] uart_s1_readdata;
  wire    [ 15: 0] uart_s1_readdata_from_sa;
  wire             uart_s1_readyfordata;
  wire             uart_s1_readyfordata_from_sa;
  wire             uart_s1_reset_n;
  wire             uart_s1_write_n;
  wire    [ 15: 0] uart_s1_writedata;
  button_pio_s1_arbitrator the_button_pio_s1
    (
      .button_pio_s1_address                           (button_pio_s1_address),
      .button_pio_s1_chipselect                        (button_pio_s1_chipselect),
      .button_pio_s1_irq                               (button_pio_s1_irq),
      .button_pio_s1_irq_from_sa                       (button_pio_s1_irq_from_sa),
      .button_pio_s1_readdata                          (button_pio_s1_readdata),
      .button_pio_s1_readdata_from_sa                  (button_pio_s1_readdata_from_sa),
      .button_pio_s1_reset_n                           (button_pio_s1_reset_n),
      .button_pio_s1_write_n                           (button_pio_s1_write_n),
      .button_pio_s1_writedata                         (button_pio_s1_writedata),
      .clk                                             (ddr3_top_phy_clk_out),
      .d1_button_pio_s1_end_xfer                       (d1_button_pio_s1_end_xfer),
      .pb_cpu_to_io_m1_address_to_slave                (pb_cpu_to_io_m1_address_to_slave),
      .pb_cpu_to_io_m1_burstcount                      (pb_cpu_to_io_m1_burstcount),
      .pb_cpu_to_io_m1_chipselect                      (pb_cpu_to_io_m1_chipselect),
      .pb_cpu_to_io_m1_granted_button_pio_s1           (pb_cpu_to_io_m1_granted_button_pio_s1),
      .pb_cpu_to_io_m1_latency_counter                 (pb_cpu_to_io_m1_latency_counter),
      .pb_cpu_to_io_m1_qualified_request_button_pio_s1 (pb_cpu_to_io_m1_qualified_request_button_pio_s1),
      .pb_cpu_to_io_m1_read                            (pb_cpu_to_io_m1_read),
      .pb_cpu_to_io_m1_read_data_valid_button_pio_s1   (pb_cpu_to_io_m1_read_data_valid_button_pio_s1),
      .pb_cpu_to_io_m1_requests_button_pio_s1          (pb_cpu_to_io_m1_requests_button_pio_s1),
      .pb_cpu_to_io_m1_write                           (pb_cpu_to_io_m1_write),
      .pb_cpu_to_io_m1_writedata                       (pb_cpu_to_io_m1_writedata),
      .reset_n                                         (ddr3_top_phy_clk_out_reset_n)
    );

  button_pio the_button_pio
    (
      .address    (button_pio_s1_address),
      .chipselect (button_pio_s1_chipselect),
      .clk        (ddr3_top_phy_clk_out),
      .in_port    (in_port_to_the_button_pio),
      .irq        (button_pio_s1_irq),
      .readdata   (button_pio_s1_readdata),
      .reset_n    (button_pio_s1_reset_n),
      .write_n    (button_pio_s1_write_n),
      .writedata  (button_pio_s1_writedata)
    );

  cpu_jtag_debug_module_arbitrator the_cpu_jtag_debug_module
    (
      .clk                                                                         (ddr3_top_phy_clk_out),
      .cpu_data_master_address_to_slave                                            (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                  (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                                 (cpu_data_master_debugaccess),
      .cpu_data_master_granted_cpu_jtag_debug_module                               (cpu_data_master_granted_cpu_jtag_debug_module),
      .cpu_data_master_latency_counter                                             (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_cpu_jtag_debug_module                     (cpu_data_master_qualified_request_cpu_jtag_debug_module),
      .cpu_data_master_read                                                        (cpu_data_master_read),
      .cpu_data_master_read_data_valid_cpu_jtag_debug_module                       (cpu_data_master_read_data_valid_cpu_jtag_debug_module),
      .cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register        (cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register),
      .cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register             (cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register),
      .cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register              (cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register),
      .cpu_data_master_requests_cpu_jtag_debug_module                              (cpu_data_master_requests_cpu_jtag_debug_module),
      .cpu_data_master_write                                                       (cpu_data_master_write),
      .cpu_data_master_writedata                                                   (cpu_data_master_writedata),
      .cpu_instruction_master_address_to_slave                                     (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_granted_cpu_jtag_debug_module                        (cpu_instruction_master_granted_cpu_jtag_debug_module),
      .cpu_instruction_master_latency_counter                                      (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_cpu_jtag_debug_module              (cpu_instruction_master_qualified_request_cpu_jtag_debug_module),
      .cpu_instruction_master_read                                                 (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_cpu_jtag_debug_module                (cpu_instruction_master_read_data_valid_cpu_jtag_debug_module),
      .cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register (cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register),
      .cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register      (cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register),
      .cpu_instruction_master_requests_cpu_jtag_debug_module                       (cpu_instruction_master_requests_cpu_jtag_debug_module),
      .cpu_jtag_debug_module_address                                               (cpu_jtag_debug_module_address),
      .cpu_jtag_debug_module_begintransfer                                         (cpu_jtag_debug_module_begintransfer),
      .cpu_jtag_debug_module_byteenable                                            (cpu_jtag_debug_module_byteenable),
      .cpu_jtag_debug_module_chipselect                                            (cpu_jtag_debug_module_chipselect),
      .cpu_jtag_debug_module_debugaccess                                           (cpu_jtag_debug_module_debugaccess),
      .cpu_jtag_debug_module_readdata                                              (cpu_jtag_debug_module_readdata),
      .cpu_jtag_debug_module_readdata_from_sa                                      (cpu_jtag_debug_module_readdata_from_sa),
      .cpu_jtag_debug_module_reset_n                                               (cpu_jtag_debug_module_reset_n),
      .cpu_jtag_debug_module_resetrequest                                          (cpu_jtag_debug_module_resetrequest),
      .cpu_jtag_debug_module_resetrequest_from_sa                                  (cpu_jtag_debug_module_resetrequest_from_sa),
      .cpu_jtag_debug_module_write                                                 (cpu_jtag_debug_module_write),
      .cpu_jtag_debug_module_writedata                                             (cpu_jtag_debug_module_writedata),
      .d1_cpu_jtag_debug_module_end_xfer                                           (d1_cpu_jtag_debug_module_end_xfer),
      .reset_n                                                                     (ddr3_top_phy_clk_out_reset_n)
    );

  cpu_data_master_arbitrator the_cpu_data_master
    (
      .button_pio_s1_irq_from_sa                                            (button_pio_s1_irq_from_sa),
      .clk                                                                  (ddr3_top_phy_clk_out),
      .cpu_data_master_address                                              (cpu_data_master_address),
      .cpu_data_master_address_to_slave                                     (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                           (cpu_data_master_byteenable),
      .cpu_data_master_granted_cpu_jtag_debug_module                        (cpu_data_master_granted_cpu_jtag_debug_module),
      .cpu_data_master_granted_pb_cpu_to_ddr3_top_s1                        (cpu_data_master_granted_pb_cpu_to_ddr3_top_s1),
      .cpu_data_master_granted_pb_cpu_to_fsm_s1                             (cpu_data_master_granted_pb_cpu_to_fsm_s1),
      .cpu_data_master_granted_pb_cpu_to_io_s1                              (cpu_data_master_granted_pb_cpu_to_io_s1),
      .cpu_data_master_irq                                                  (cpu_data_master_irq),
      .cpu_data_master_latency_counter                                      (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_cpu_jtag_debug_module              (cpu_data_master_qualified_request_cpu_jtag_debug_module),
      .cpu_data_master_qualified_request_pb_cpu_to_ddr3_top_s1              (cpu_data_master_qualified_request_pb_cpu_to_ddr3_top_s1),
      .cpu_data_master_qualified_request_pb_cpu_to_fsm_s1                   (cpu_data_master_qualified_request_pb_cpu_to_fsm_s1),
      .cpu_data_master_qualified_request_pb_cpu_to_io_s1                    (cpu_data_master_qualified_request_pb_cpu_to_io_s1),
      .cpu_data_master_read                                                 (cpu_data_master_read),
      .cpu_data_master_read_data_valid_cpu_jtag_debug_module                (cpu_data_master_read_data_valid_cpu_jtag_debug_module),
      .cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1                (cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1),
      .cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register (cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register),
      .cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1                     (cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1),
      .cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register      (cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register),
      .cpu_data_master_read_data_valid_pb_cpu_to_io_s1                      (cpu_data_master_read_data_valid_pb_cpu_to_io_s1),
      .cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register       (cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register),
      .cpu_data_master_readdata                                             (cpu_data_master_readdata),
      .cpu_data_master_readdatavalid                                        (cpu_data_master_readdatavalid),
      .cpu_data_master_requests_cpu_jtag_debug_module                       (cpu_data_master_requests_cpu_jtag_debug_module),
      .cpu_data_master_requests_pb_cpu_to_ddr3_top_s1                       (cpu_data_master_requests_pb_cpu_to_ddr3_top_s1),
      .cpu_data_master_requests_pb_cpu_to_fsm_s1                            (cpu_data_master_requests_pb_cpu_to_fsm_s1),
      .cpu_data_master_requests_pb_cpu_to_io_s1                             (cpu_data_master_requests_pb_cpu_to_io_s1),
      .cpu_data_master_waitrequest                                          (cpu_data_master_waitrequest),
      .cpu_data_master_write                                                (cpu_data_master_write),
      .cpu_data_master_writedata                                            (cpu_data_master_writedata),
      .cpu_jtag_debug_module_readdata_from_sa                               (cpu_jtag_debug_module_readdata_from_sa),
      .d1_cpu_jtag_debug_module_end_xfer                                    (d1_cpu_jtag_debug_module_end_xfer),
      .d1_pb_cpu_to_ddr3_top_s1_end_xfer                                    (d1_pb_cpu_to_ddr3_top_s1_end_xfer),
      .d1_pb_cpu_to_fsm_s1_end_xfer                                         (d1_pb_cpu_to_fsm_s1_end_xfer),
      .d1_pb_cpu_to_io_s1_end_xfer                                          (d1_pb_cpu_to_io_s1_end_xfer),
      .dipsw_pio_s1_irq_from_sa                                             (dipsw_pio_s1_irq_from_sa),
      .jtag_uart_avalon_jtag_slave_irq_from_sa                              (jtag_uart_avalon_jtag_slave_irq_from_sa),
      .pb_cpu_to_ddr3_top_s1_readdata_from_sa                               (pb_cpu_to_ddr3_top_s1_readdata_from_sa),
      .pb_cpu_to_ddr3_top_s1_waitrequest_from_sa                            (pb_cpu_to_ddr3_top_s1_waitrequest_from_sa),
      .pb_cpu_to_fsm_s1_readdata_from_sa                                    (pb_cpu_to_fsm_s1_readdata_from_sa),
      .pb_cpu_to_fsm_s1_waitrequest_from_sa                                 (pb_cpu_to_fsm_s1_waitrequest_from_sa),
      .pb_cpu_to_io_s1_readdata_from_sa                                     (pb_cpu_to_io_s1_readdata_from_sa),
      .pb_cpu_to_io_s1_waitrequest_from_sa                                  (pb_cpu_to_io_s1_waitrequest_from_sa),
      .reset_n                                                              (ddr3_top_phy_clk_out_reset_n),
      .sgdma_rx_csr_irq_from_sa                                             (sgdma_rx_csr_irq_from_sa),
      .sgdma_tx_csr_irq_from_sa                                             (sgdma_tx_csr_irq_from_sa),
      .timer_1ms_s1_irq_from_sa                                             (timer_1ms_s1_irq_from_sa),
      .uart_s1_irq_from_sa                                                  (uart_s1_irq_from_sa)
    );

  cpu_instruction_master_arbitrator the_cpu_instruction_master
    (
      .clk                                                                         (ddr3_top_phy_clk_out),
      .cpu_instruction_master_address                                              (cpu_instruction_master_address),
      .cpu_instruction_master_address_to_slave                                     (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_granted_cpu_jtag_debug_module                        (cpu_instruction_master_granted_cpu_jtag_debug_module),
      .cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1                        (cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1),
      .cpu_instruction_master_granted_pb_cpu_to_fsm_s1                             (cpu_instruction_master_granted_pb_cpu_to_fsm_s1),
      .cpu_instruction_master_latency_counter                                      (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_cpu_jtag_debug_module              (cpu_instruction_master_qualified_request_cpu_jtag_debug_module),
      .cpu_instruction_master_qualified_request_pb_cpu_to_ddr3_top_s1              (cpu_instruction_master_qualified_request_pb_cpu_to_ddr3_top_s1),
      .cpu_instruction_master_qualified_request_pb_cpu_to_fsm_s1                   (cpu_instruction_master_qualified_request_pb_cpu_to_fsm_s1),
      .cpu_instruction_master_read                                                 (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_cpu_jtag_debug_module                (cpu_instruction_master_read_data_valid_cpu_jtag_debug_module),
      .cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1                (cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1),
      .cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register (cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register),
      .cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1                     (cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1),
      .cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register      (cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register),
      .cpu_instruction_master_readdata                                             (cpu_instruction_master_readdata),
      .cpu_instruction_master_readdatavalid                                        (cpu_instruction_master_readdatavalid),
      .cpu_instruction_master_requests_cpu_jtag_debug_module                       (cpu_instruction_master_requests_cpu_jtag_debug_module),
      .cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1                       (cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1),
      .cpu_instruction_master_requests_pb_cpu_to_fsm_s1                            (cpu_instruction_master_requests_pb_cpu_to_fsm_s1),
      .cpu_instruction_master_waitrequest                                          (cpu_instruction_master_waitrequest),
      .cpu_jtag_debug_module_readdata_from_sa                                      (cpu_jtag_debug_module_readdata_from_sa),
      .d1_cpu_jtag_debug_module_end_xfer                                           (d1_cpu_jtag_debug_module_end_xfer),
      .d1_pb_cpu_to_ddr3_top_s1_end_xfer                                           (d1_pb_cpu_to_ddr3_top_s1_end_xfer),
      .d1_pb_cpu_to_fsm_s1_end_xfer                                                (d1_pb_cpu_to_fsm_s1_end_xfer),
      .pb_cpu_to_ddr3_top_s1_readdata_from_sa                                      (pb_cpu_to_ddr3_top_s1_readdata_from_sa),
      .pb_cpu_to_ddr3_top_s1_waitrequest_from_sa                                   (pb_cpu_to_ddr3_top_s1_waitrequest_from_sa),
      .pb_cpu_to_fsm_s1_readdata_from_sa                                           (pb_cpu_to_fsm_s1_readdata_from_sa),
      .pb_cpu_to_fsm_s1_waitrequest_from_sa                                        (pb_cpu_to_fsm_s1_waitrequest_from_sa),
      .reset_n                                                                     (ddr3_top_phy_clk_out_reset_n)
    );

  cpu_tightly_coupled_data_master_0_arbitrator the_cpu_tightly_coupled_data_master_0
    (
      .clk                                                                    (ddr3_top_phy_clk_out),
      .cpu_tightly_coupled_data_master_0_address                              (cpu_tightly_coupled_data_master_0_address),
      .cpu_tightly_coupled_data_master_0_address_to_slave                     (cpu_tightly_coupled_data_master_0_address_to_slave),
      .cpu_tightly_coupled_data_master_0_byteenable                           (cpu_tightly_coupled_data_master_0_byteenable),
      .cpu_tightly_coupled_data_master_0_clken                                (cpu_tightly_coupled_data_master_0_clken),
      .cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2           (cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2),
      .cpu_tightly_coupled_data_master_0_latency_counter                      (cpu_tightly_coupled_data_master_0_latency_counter),
      .cpu_tightly_coupled_data_master_0_qualified_request_tlb_miss_ram_1k_s2 (cpu_tightly_coupled_data_master_0_qualified_request_tlb_miss_ram_1k_s2),
      .cpu_tightly_coupled_data_master_0_read                                 (cpu_tightly_coupled_data_master_0_read),
      .cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2   (cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2),
      .cpu_tightly_coupled_data_master_0_readdata                             (cpu_tightly_coupled_data_master_0_readdata),
      .cpu_tightly_coupled_data_master_0_readdatavalid                        (cpu_tightly_coupled_data_master_0_readdatavalid),
      .cpu_tightly_coupled_data_master_0_requests_tlb_miss_ram_1k_s2          (cpu_tightly_coupled_data_master_0_requests_tlb_miss_ram_1k_s2),
      .cpu_tightly_coupled_data_master_0_waitrequest                          (cpu_tightly_coupled_data_master_0_waitrequest),
      .cpu_tightly_coupled_data_master_0_write                                (cpu_tightly_coupled_data_master_0_write),
      .cpu_tightly_coupled_data_master_0_writedata                            (cpu_tightly_coupled_data_master_0_writedata),
      .d1_tlb_miss_ram_1k_s2_end_xfer                                         (d1_tlb_miss_ram_1k_s2_end_xfer),
      .reset_n                                                                (ddr3_top_phy_clk_out_reset_n),
      .tlb_miss_ram_1k_s2_readdata_from_sa                                    (tlb_miss_ram_1k_s2_readdata_from_sa)
    );

  cpu_tightly_coupled_instruction_master_0_arbitrator the_cpu_tightly_coupled_instruction_master_0
    (
      .clk                                                                           (ddr3_top_phy_clk_out),
      .cpu_tightly_coupled_instruction_master_0_address                              (cpu_tightly_coupled_instruction_master_0_address),
      .cpu_tightly_coupled_instruction_master_0_address_to_slave                     (cpu_tightly_coupled_instruction_master_0_address_to_slave),
      .cpu_tightly_coupled_instruction_master_0_clken                                (cpu_tightly_coupled_instruction_master_0_clken),
      .cpu_tightly_coupled_instruction_master_0_granted_tlb_miss_ram_1k_s1           (cpu_tightly_coupled_instruction_master_0_granted_tlb_miss_ram_1k_s1),
      .cpu_tightly_coupled_instruction_master_0_latency_counter                      (cpu_tightly_coupled_instruction_master_0_latency_counter),
      .cpu_tightly_coupled_instruction_master_0_qualified_request_tlb_miss_ram_1k_s1 (cpu_tightly_coupled_instruction_master_0_qualified_request_tlb_miss_ram_1k_s1),
      .cpu_tightly_coupled_instruction_master_0_read                                 (cpu_tightly_coupled_instruction_master_0_read),
      .cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1   (cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1),
      .cpu_tightly_coupled_instruction_master_0_readdata                             (cpu_tightly_coupled_instruction_master_0_readdata),
      .cpu_tightly_coupled_instruction_master_0_readdatavalid                        (cpu_tightly_coupled_instruction_master_0_readdatavalid),
      .cpu_tightly_coupled_instruction_master_0_requests_tlb_miss_ram_1k_s1          (cpu_tightly_coupled_instruction_master_0_requests_tlb_miss_ram_1k_s1),
      .cpu_tightly_coupled_instruction_master_0_waitrequest                          (cpu_tightly_coupled_instruction_master_0_waitrequest),
      .d1_tlb_miss_ram_1k_s1_end_xfer                                                (d1_tlb_miss_ram_1k_s1_end_xfer),
      .reset_n                                                                       (ddr3_top_phy_clk_out_reset_n),
      .tlb_miss_ram_1k_s1_readdata_from_sa                                           (tlb_miss_ram_1k_s1_readdata_from_sa)
    );

  cpu the_cpu
    (
      .clk                                   (ddr3_top_phy_clk_out),
      .d_address                             (cpu_data_master_address),
      .d_byteenable                          (cpu_data_master_byteenable),
      .d_irq                                 (cpu_data_master_irq),
      .d_read                                (cpu_data_master_read),
      .d_readdata                            (cpu_data_master_readdata),
      .d_readdatavalid                       (cpu_data_master_readdatavalid),
      .d_waitrequest                         (cpu_data_master_waitrequest),
      .d_write                               (cpu_data_master_write),
      .d_writedata                           (cpu_data_master_writedata),
      .dcm0_address                          (cpu_tightly_coupled_data_master_0_address),
      .dcm0_byteenable                       (cpu_tightly_coupled_data_master_0_byteenable),
      .dcm0_clken                            (cpu_tightly_coupled_data_master_0_clken),
      .dcm0_read                             (cpu_tightly_coupled_data_master_0_read),
      .dcm0_readdata                         (cpu_tightly_coupled_data_master_0_readdata),
      .dcm0_readdatavalid                    (cpu_tightly_coupled_data_master_0_readdatavalid),
      .dcm0_waitrequest                      (cpu_tightly_coupled_data_master_0_waitrequest),
      .dcm0_write                            (cpu_tightly_coupled_data_master_0_write),
      .dcm0_writedata                        (cpu_tightly_coupled_data_master_0_writedata),
      .i_address                             (cpu_instruction_master_address),
      .i_read                                (cpu_instruction_master_read),
      .i_readdata                            (cpu_instruction_master_readdata),
      .i_readdatavalid                       (cpu_instruction_master_readdatavalid),
      .i_waitrequest                         (cpu_instruction_master_waitrequest),
      .icm0_address                          (cpu_tightly_coupled_instruction_master_0_address),
      .icm0_clken                            (cpu_tightly_coupled_instruction_master_0_clken),
      .icm0_read                             (cpu_tightly_coupled_instruction_master_0_read),
      .icm0_readdata                         (cpu_tightly_coupled_instruction_master_0_readdata),
      .icm0_readdatavalid                    (cpu_tightly_coupled_instruction_master_0_readdatavalid),
      .icm0_waitrequest                      (cpu_tightly_coupled_instruction_master_0_waitrequest),
      .jtag_debug_module_address             (cpu_jtag_debug_module_address),
      .jtag_debug_module_begintransfer       (cpu_jtag_debug_module_begintransfer),
      .jtag_debug_module_byteenable          (cpu_jtag_debug_module_byteenable),
      .jtag_debug_module_debugaccess         (cpu_jtag_debug_module_debugaccess),
      .jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),
      .jtag_debug_module_readdata            (cpu_jtag_debug_module_readdata),
      .jtag_debug_module_resetrequest        (cpu_jtag_debug_module_resetrequest),
      .jtag_debug_module_select              (cpu_jtag_debug_module_chipselect),
      .jtag_debug_module_write               (cpu_jtag_debug_module_write),
      .jtag_debug_module_writedata           (cpu_jtag_debug_module_writedata),
      .reset_n                               (cpu_jtag_debug_module_reset_n)
    );

  ddr3_top_s1_arbitrator the_ddr3_top_s1
    (
      .clk                                                              (ddr3_top_phy_clk_out),
      .d1_ddr3_top_s1_end_xfer                                          (d1_ddr3_top_s1_end_xfer),
      .ddr3_top_s1_address                                              (ddr3_top_s1_address),
      .ddr3_top_s1_beginbursttransfer                                   (ddr3_top_s1_beginbursttransfer),
      .ddr3_top_s1_burstcount                                           (ddr3_top_s1_burstcount),
      .ddr3_top_s1_byteenable                                           (ddr3_top_s1_byteenable),
      .ddr3_top_s1_read                                                 (ddr3_top_s1_read),
      .ddr3_top_s1_readdata                                             (ddr3_top_s1_readdata),
      .ddr3_top_s1_readdata_from_sa                                     (ddr3_top_s1_readdata_from_sa),
      .ddr3_top_s1_readdatavalid                                        (ddr3_top_s1_readdatavalid),
      .ddr3_top_s1_resetrequest_n                                       (ddr3_top_s1_resetrequest_n),
      .ddr3_top_s1_resetrequest_n_from_sa                               (ddr3_top_s1_resetrequest_n_from_sa),
      .ddr3_top_s1_waitrequest_n                                        (ddr3_top_s1_waitrequest_n),
      .ddr3_top_s1_waitrequest_n_from_sa                                (ddr3_top_s1_waitrequest_n_from_sa),
      .ddr3_top_s1_write                                                (ddr3_top_s1_write),
      .ddr3_top_s1_writedata                                            (ddr3_top_s1_writedata),
      .pb_cpu_to_ddr3_top_m1_address_to_slave                           (pb_cpu_to_ddr3_top_m1_address_to_slave),
      .pb_cpu_to_ddr3_top_m1_burstcount                                 (pb_cpu_to_ddr3_top_m1_burstcount),
      .pb_cpu_to_ddr3_top_m1_byteenable                                 (pb_cpu_to_ddr3_top_m1_byteenable),
      .pb_cpu_to_ddr3_top_m1_chipselect                                 (pb_cpu_to_ddr3_top_m1_chipselect),
      .pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1                        (pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1),
      .pb_cpu_to_ddr3_top_m1_latency_counter                            (pb_cpu_to_ddr3_top_m1_latency_counter),
      .pb_cpu_to_ddr3_top_m1_qualified_request_ddr3_top_s1              (pb_cpu_to_ddr3_top_m1_qualified_request_ddr3_top_s1),
      .pb_cpu_to_ddr3_top_m1_read                                       (pb_cpu_to_ddr3_top_m1_read),
      .pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1                (pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1),
      .pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register (pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register),
      .pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1                       (pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1),
      .pb_cpu_to_ddr3_top_m1_write                                      (pb_cpu_to_ddr3_top_m1_write),
      .pb_cpu_to_ddr3_top_m1_writedata                                  (pb_cpu_to_ddr3_top_m1_writedata),
      .pb_dma_to_ddr3_top_m1_address_to_slave                           (pb_dma_to_ddr3_top_m1_address_to_slave),
      .pb_dma_to_ddr3_top_m1_burstcount                                 (pb_dma_to_ddr3_top_m1_burstcount),
      .pb_dma_to_ddr3_top_m1_byteenable                                 (pb_dma_to_ddr3_top_m1_byteenable),
      .pb_dma_to_ddr3_top_m1_chipselect                                 (pb_dma_to_ddr3_top_m1_chipselect),
      .pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1                        (pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1),
      .pb_dma_to_ddr3_top_m1_latency_counter                            (pb_dma_to_ddr3_top_m1_latency_counter),
      .pb_dma_to_ddr3_top_m1_qualified_request_ddr3_top_s1              (pb_dma_to_ddr3_top_m1_qualified_request_ddr3_top_s1),
      .pb_dma_to_ddr3_top_m1_read                                       (pb_dma_to_ddr3_top_m1_read),
      .pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1                (pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1),
      .pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register (pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register),
      .pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1                       (pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1),
      .pb_dma_to_ddr3_top_m1_write                                      (pb_dma_to_ddr3_top_m1_write),
      .pb_dma_to_ddr3_top_m1_writedata                                  (pb_dma_to_ddr3_top_m1_writedata),
      .reset_n                                                          (ddr3_top_phy_clk_out_reset_n)
    );

  //ddr3_top_aux_full_rate_clk_out out_clk assignment, which is an e_assign
  assign ddr3_top_aux_full_rate_clk_out = out_clk_ddr3_top_aux_full_rate_clk;

  //ddr3_top_aux_half_rate_clk_out out_clk assignment, which is an e_assign
  assign ddr3_top_aux_half_rate_clk_out = out_clk_ddr3_top_aux_half_rate_clk;

  //ddr3_top_phy_clk_out out_clk assignment, which is an e_assign
  assign ddr3_top_phy_clk_out = out_clk_ddr3_top_phy_clk;

  //reset is asserted asynchronously and deasserted synchronously
  ghrd_4sgx230_sopc_reset_clkin_100_domain_synch_module ghrd_4sgx230_sopc_reset_clkin_100_domain_synch
    (
      .clk      (clkin_100),
      .data_in  (1'b1),
      .data_out (clkin_100_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset sources mux, which is an e_mux
  assign reset_n_sources = ~(~reset_n |
    0 |
    0 |
    cpu_jtag_debug_module_resetrequest_from_sa |
    cpu_jtag_debug_module_resetrequest_from_sa |
    ~ddr3_top_s1_resetrequest_n_from_sa |
    ~ddr3_top_s1_resetrequest_n_from_sa);

  ddr3_top the_ddr3_top
    (
      .aux_full_rate_clk     (out_clk_ddr3_top_aux_full_rate_clk),
      .aux_half_rate_clk     (out_clk_ddr3_top_aux_half_rate_clk),
      .aux_scan_clk          (aux_scan_clk_from_the_ddr3_top),
      .aux_scan_clk_reset_n  (aux_scan_clk_reset_n_from_the_ddr3_top),
      .dll_reference_clk     (dll_reference_clk_from_the_ddr3_top),
      .dqs_delay_ctrl_export (dqs_delay_ctrl_export_from_the_ddr3_top),
      .global_reset_n        (global_reset_n_to_the_ddr3_top),
      .local_address         (ddr3_top_s1_address),
      .local_be              (ddr3_top_s1_byteenable),
      .local_burstbegin      (ddr3_top_s1_beginbursttransfer),
      .local_init_done       (local_init_done_from_the_ddr3_top),
      .local_rdata           (ddr3_top_s1_readdata),
      .local_rdata_valid     (ddr3_top_s1_readdatavalid),
      .local_read_req        (ddr3_top_s1_read),
      .local_ready           (ddr3_top_s1_waitrequest_n),
      .local_refresh_ack     (local_refresh_ack_from_the_ddr3_top),
      .local_size            (ddr3_top_s1_burstcount),
      .local_wdata           (ddr3_top_s1_writedata),
      .local_wdata_req       (local_wdata_req_from_the_ddr3_top),
      .local_write_req       (ddr3_top_s1_write),
      .mem_addr              (mem_addr_from_the_ddr3_top),
      .mem_ba                (mem_ba_from_the_ddr3_top),
      .mem_cas_n             (mem_cas_n_from_the_ddr3_top),
      .mem_cke               (mem_cke_from_the_ddr3_top),
      .mem_clk               (mem_clk_to_and_from_the_ddr3_top),
      .mem_clk_n             (mem_clk_n_to_and_from_the_ddr3_top),
      .mem_cs_n              (mem_cs_n_from_the_ddr3_top),
      .mem_dm                (mem_dm_from_the_ddr3_top),
      .mem_dq                (mem_dq_to_and_from_the_ddr3_top),
      .mem_dqs               (mem_dqs_to_and_from_the_ddr3_top),
      .mem_dqsn              (mem_dqsn_to_and_from_the_ddr3_top),
      .mem_odt               (mem_odt_from_the_ddr3_top),
      .mem_ras_n             (mem_ras_n_from_the_ddr3_top),
      .mem_reset_n           (mem_reset_n_from_the_ddr3_top),
      .mem_we_n              (mem_we_n_from_the_ddr3_top),
      .oct_ctl_rs_value      (oct_ctl_rs_value_to_the_ddr3_top),
      .oct_ctl_rt_value      (oct_ctl_rt_value_to_the_ddr3_top),
      .phy_clk               (out_clk_ddr3_top_phy_clk),
      .pll_ref_clk           (clkin_100),
      .reset_phy_clk_n       (reset_phy_clk_n_from_the_ddr3_top),
      .reset_request_n       (ddr3_top_s1_resetrequest_n),
      .soft_reset_n          (clkin_100_reset_n)
    );

  descriptor_memory_s1_arbitrator the_descriptor_memory_s1
    (
      .clk                                                                   (ddr3_top_phy_clk_out),
      .d1_descriptor_memory_s1_end_xfer                                      (d1_descriptor_memory_s1_end_xfer),
      .descriptor_memory_s1_address                                          (descriptor_memory_s1_address),
      .descriptor_memory_s1_byteenable                                       (descriptor_memory_s1_byteenable),
      .descriptor_memory_s1_chipselect                                       (descriptor_memory_s1_chipselect),
      .descriptor_memory_s1_clken                                            (descriptor_memory_s1_clken),
      .descriptor_memory_s1_readdata                                         (descriptor_memory_s1_readdata),
      .descriptor_memory_s1_readdata_from_sa                                 (descriptor_memory_s1_readdata_from_sa),
      .descriptor_memory_s1_reset                                            (descriptor_memory_s1_reset),
      .descriptor_memory_s1_write                                            (descriptor_memory_s1_write),
      .descriptor_memory_s1_writedata                                        (descriptor_memory_s1_writedata),
      .pb_cpu_to_io_m1_address_to_slave                                      (pb_cpu_to_io_m1_address_to_slave),
      .pb_cpu_to_io_m1_burstcount                                            (pb_cpu_to_io_m1_burstcount),
      .pb_cpu_to_io_m1_byteenable                                            (pb_cpu_to_io_m1_byteenable),
      .pb_cpu_to_io_m1_chipselect                                            (pb_cpu_to_io_m1_chipselect),
      .pb_cpu_to_io_m1_granted_descriptor_memory_s1                          (pb_cpu_to_io_m1_granted_descriptor_memory_s1),
      .pb_cpu_to_io_m1_latency_counter                                       (pb_cpu_to_io_m1_latency_counter),
      .pb_cpu_to_io_m1_qualified_request_descriptor_memory_s1                (pb_cpu_to_io_m1_qualified_request_descriptor_memory_s1),
      .pb_cpu_to_io_m1_read                                                  (pb_cpu_to_io_m1_read),
      .pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1                  (pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1),
      .pb_cpu_to_io_m1_requests_descriptor_memory_s1                         (pb_cpu_to_io_m1_requests_descriptor_memory_s1),
      .pb_cpu_to_io_m1_write                                                 (pb_cpu_to_io_m1_write),
      .pb_cpu_to_io_m1_writedata                                             (pb_cpu_to_io_m1_writedata),
      .pb_dma_to_descriptor_memory_m1_address_to_slave                       (pb_dma_to_descriptor_memory_m1_address_to_slave),
      .pb_dma_to_descriptor_memory_m1_burstcount                             (pb_dma_to_descriptor_memory_m1_burstcount),
      .pb_dma_to_descriptor_memory_m1_byteenable                             (pb_dma_to_descriptor_memory_m1_byteenable),
      .pb_dma_to_descriptor_memory_m1_chipselect                             (pb_dma_to_descriptor_memory_m1_chipselect),
      .pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1           (pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1),
      .pb_dma_to_descriptor_memory_m1_latency_counter                        (pb_dma_to_descriptor_memory_m1_latency_counter),
      .pb_dma_to_descriptor_memory_m1_qualified_request_descriptor_memory_s1 (pb_dma_to_descriptor_memory_m1_qualified_request_descriptor_memory_s1),
      .pb_dma_to_descriptor_memory_m1_read                                   (pb_dma_to_descriptor_memory_m1_read),
      .pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1   (pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1),
      .pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1          (pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1),
      .pb_dma_to_descriptor_memory_m1_write                                  (pb_dma_to_descriptor_memory_m1_write),
      .pb_dma_to_descriptor_memory_m1_writedata                              (pb_dma_to_descriptor_memory_m1_writedata),
      .reset_n                                                               (ddr3_top_phy_clk_out_reset_n)
    );

  descriptor_memory the_descriptor_memory
    (
      .address    (descriptor_memory_s1_address),
      .byteenable (descriptor_memory_s1_byteenable),
      .chipselect (descriptor_memory_s1_chipselect),
      .clk        (ddr3_top_phy_clk_out),
      .clken      (descriptor_memory_s1_clken),
      .readdata   (descriptor_memory_s1_readdata),
      .reset      (descriptor_memory_s1_reset),
      .write      (descriptor_memory_s1_write),
      .writedata  (descriptor_memory_s1_writedata)
    );

  dipsw_pio_s1_arbitrator the_dipsw_pio_s1
    (
      .clk                                            (ddr3_top_phy_clk_out),
      .d1_dipsw_pio_s1_end_xfer                       (d1_dipsw_pio_s1_end_xfer),
      .dipsw_pio_s1_address                           (dipsw_pio_s1_address),
      .dipsw_pio_s1_chipselect                        (dipsw_pio_s1_chipselect),
      .dipsw_pio_s1_irq                               (dipsw_pio_s1_irq),
      .dipsw_pio_s1_irq_from_sa                       (dipsw_pio_s1_irq_from_sa),
      .dipsw_pio_s1_readdata                          (dipsw_pio_s1_readdata),
      .dipsw_pio_s1_readdata_from_sa                  (dipsw_pio_s1_readdata_from_sa),
      .dipsw_pio_s1_reset_n                           (dipsw_pio_s1_reset_n),
      .dipsw_pio_s1_write_n                           (dipsw_pio_s1_write_n),
      .dipsw_pio_s1_writedata                         (dipsw_pio_s1_writedata),
      .pb_cpu_to_io_m1_address_to_slave               (pb_cpu_to_io_m1_address_to_slave),
      .pb_cpu_to_io_m1_burstcount                     (pb_cpu_to_io_m1_burstcount),
      .pb_cpu_to_io_m1_byteenable                     (pb_cpu_to_io_m1_byteenable),
      .pb_cpu_to_io_m1_chipselect                     (pb_cpu_to_io_m1_chipselect),
      .pb_cpu_to_io_m1_granted_dipsw_pio_s1           (pb_cpu_to_io_m1_granted_dipsw_pio_s1),
      .pb_cpu_to_io_m1_latency_counter                (pb_cpu_to_io_m1_latency_counter),
      .pb_cpu_to_io_m1_qualified_request_dipsw_pio_s1 (pb_cpu_to_io_m1_qualified_request_dipsw_pio_s1),
      .pb_cpu_to_io_m1_read                           (pb_cpu_to_io_m1_read),
      .pb_cpu_to_io_m1_read_data_valid_dipsw_pio_s1   (pb_cpu_to_io_m1_read_data_valid_dipsw_pio_s1),
      .pb_cpu_to_io_m1_requests_dipsw_pio_s1          (pb_cpu_to_io_m1_requests_dipsw_pio_s1),
      .pb_cpu_to_io_m1_write                          (pb_cpu_to_io_m1_write),
      .pb_cpu_to_io_m1_writedata                      (pb_cpu_to_io_m1_writedata),
      .reset_n                                        (ddr3_top_phy_clk_out_reset_n)
    );

  dipsw_pio the_dipsw_pio
    (
      .address    (dipsw_pio_s1_address),
      .chipselect (dipsw_pio_s1_chipselect),
      .clk        (ddr3_top_phy_clk_out),
      .in_port    (in_port_to_the_dipsw_pio),
      .irq        (dipsw_pio_s1_irq),
      .readdata   (dipsw_pio_s1_readdata),
      .reset_n    (dipsw_pio_s1_reset_n),
      .write_n    (dipsw_pio_s1_write_n),
      .writedata  (dipsw_pio_s1_writedata)
    );

  jtag_uart_avalon_jtag_slave_arbitrator the_jtag_uart_avalon_jtag_slave
    (
      .clk                                                           (ddr3_top_phy_clk_out),
      .d1_jtag_uart_avalon_jtag_slave_end_xfer                       (d1_jtag_uart_avalon_jtag_slave_end_xfer),
      .jtag_uart_avalon_jtag_slave_address                           (jtag_uart_avalon_jtag_slave_address),
      .jtag_uart_avalon_jtag_slave_chipselect                        (jtag_uart_avalon_jtag_slave_chipselect),
      .jtag_uart_avalon_jtag_slave_dataavailable                     (jtag_uart_avalon_jtag_slave_dataavailable),
      .jtag_uart_avalon_jtag_slave_dataavailable_from_sa             (jtag_uart_avalon_jtag_slave_dataavailable_from_sa),
      .jtag_uart_avalon_jtag_slave_irq                               (jtag_uart_avalon_jtag_slave_irq),
      .jtag_uart_avalon_jtag_slave_irq_from_sa                       (jtag_uart_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_avalon_jtag_slave_read_n                            (jtag_uart_avalon_jtag_slave_read_n),
      .jtag_uart_avalon_jtag_slave_readdata                          (jtag_uart_avalon_jtag_slave_readdata),
      .jtag_uart_avalon_jtag_slave_readdata_from_sa                  (jtag_uart_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_readyfordata                      (jtag_uart_avalon_jtag_slave_readyfordata),
      .jtag_uart_avalon_jtag_slave_readyfordata_from_sa              (jtag_uart_avalon_jtag_slave_readyfordata_from_sa),
      .jtag_uart_avalon_jtag_slave_reset_n                           (jtag_uart_avalon_jtag_slave_reset_n),
      .jtag_uart_avalon_jtag_slave_waitrequest                       (jtag_uart_avalon_jtag_slave_waitrequest),
      .jtag_uart_avalon_jtag_slave_waitrequest_from_sa               (jtag_uart_avalon_jtag_slave_waitrequest_from_sa),
      .jtag_uart_avalon_jtag_slave_write_n                           (jtag_uart_avalon_jtag_slave_write_n),
      .jtag_uart_avalon_jtag_slave_writedata                         (jtag_uart_avalon_jtag_slave_writedata),
      .pb_cpu_to_io_m1_address_to_slave                              (pb_cpu_to_io_m1_address_to_slave),
      .pb_cpu_to_io_m1_burstcount                                    (pb_cpu_to_io_m1_burstcount),
      .pb_cpu_to_io_m1_chipselect                                    (pb_cpu_to_io_m1_chipselect),
      .pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave           (pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave),
      .pb_cpu_to_io_m1_latency_counter                               (pb_cpu_to_io_m1_latency_counter),
      .pb_cpu_to_io_m1_qualified_request_jtag_uart_avalon_jtag_slave (pb_cpu_to_io_m1_qualified_request_jtag_uart_avalon_jtag_slave),
      .pb_cpu_to_io_m1_read                                          (pb_cpu_to_io_m1_read),
      .pb_cpu_to_io_m1_read_data_valid_jtag_uart_avalon_jtag_slave   (pb_cpu_to_io_m1_read_data_valid_jtag_uart_avalon_jtag_slave),
      .pb_cpu_to_io_m1_requests_jtag_uart_avalon_jtag_slave          (pb_cpu_to_io_m1_requests_jtag_uart_avalon_jtag_slave),
      .pb_cpu_to_io_m1_write                                         (pb_cpu_to_io_m1_write),
      .pb_cpu_to_io_m1_writedata                                     (pb_cpu_to_io_m1_writedata),
      .reset_n                                                       (ddr3_top_phy_clk_out_reset_n)
    );

  jtag_uart the_jtag_uart
    (
      .av_address     (jtag_uart_avalon_jtag_slave_address),
      .av_chipselect  (jtag_uart_avalon_jtag_slave_chipselect),
      .av_irq         (jtag_uart_avalon_jtag_slave_irq),
      .av_read_n      (jtag_uart_avalon_jtag_slave_read_n),
      .av_readdata    (jtag_uart_avalon_jtag_slave_readdata),
      .av_waitrequest (jtag_uart_avalon_jtag_slave_waitrequest),
      .av_write_n     (jtag_uart_avalon_jtag_slave_write_n),
      .av_writedata   (jtag_uart_avalon_jtag_slave_writedata),
      .clk            (ddr3_top_phy_clk_out),
      .dataavailable  (jtag_uart_avalon_jtag_slave_dataavailable),
      .readyfordata   (jtag_uart_avalon_jtag_slave_readyfordata),
      .rst_n          (jtag_uart_avalon_jtag_slave_reset_n)
    );

  led_pio_s1_arbitrator the_led_pio_s1
    (
      .clk                                          (ddr3_top_phy_clk_out),
      .d1_led_pio_s1_end_xfer                       (d1_led_pio_s1_end_xfer),
      .led_pio_s1_address                           (led_pio_s1_address),
      .led_pio_s1_chipselect                        (led_pio_s1_chipselect),
      .led_pio_s1_readdata                          (led_pio_s1_readdata),
      .led_pio_s1_readdata_from_sa                  (led_pio_s1_readdata_from_sa),
      .led_pio_s1_reset_n                           (led_pio_s1_reset_n),
      .led_pio_s1_write_n                           (led_pio_s1_write_n),
      .led_pio_s1_writedata                         (led_pio_s1_writedata),
      .pb_cpu_to_io_m1_address_to_slave             (pb_cpu_to_io_m1_address_to_slave),
      .pb_cpu_to_io_m1_burstcount                   (pb_cpu_to_io_m1_burstcount),
      .pb_cpu_to_io_m1_chipselect                   (pb_cpu_to_io_m1_chipselect),
      .pb_cpu_to_io_m1_granted_led_pio_s1           (pb_cpu_to_io_m1_granted_led_pio_s1),
      .pb_cpu_to_io_m1_latency_counter              (pb_cpu_to_io_m1_latency_counter),
      .pb_cpu_to_io_m1_qualified_request_led_pio_s1 (pb_cpu_to_io_m1_qualified_request_led_pio_s1),
      .pb_cpu_to_io_m1_read                         (pb_cpu_to_io_m1_read),
      .pb_cpu_to_io_m1_read_data_valid_led_pio_s1   (pb_cpu_to_io_m1_read_data_valid_led_pio_s1),
      .pb_cpu_to_io_m1_requests_led_pio_s1          (pb_cpu_to_io_m1_requests_led_pio_s1),
      .pb_cpu_to_io_m1_write                        (pb_cpu_to_io_m1_write),
      .pb_cpu_to_io_m1_writedata                    (pb_cpu_to_io_m1_writedata),
      .reset_n                                      (ddr3_top_phy_clk_out_reset_n)
    );

  led_pio the_led_pio
    (
      .address    (led_pio_s1_address),
      .chipselect (led_pio_s1_chipselect),
      .clk        (ddr3_top_phy_clk_out),
      .out_port   (out_port_from_the_led_pio),
      .readdata   (led_pio_s1_readdata),
      .reset_n    (led_pio_s1_reset_n),
      .write_n    (led_pio_s1_write_n),
      .writedata  (led_pio_s1_writedata)
    );

  pb_cpu_to_ddr3_top_s1_arbitrator the_pb_cpu_to_ddr3_top_s1
    (
      .clk                                                                         (ddr3_top_phy_clk_out),
      .cpu_data_master_address_to_slave                                            (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                  (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                                 (cpu_data_master_debugaccess),
      .cpu_data_master_granted_pb_cpu_to_ddr3_top_s1                               (cpu_data_master_granted_pb_cpu_to_ddr3_top_s1),
      .cpu_data_master_latency_counter                                             (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_pb_cpu_to_ddr3_top_s1                     (cpu_data_master_qualified_request_pb_cpu_to_ddr3_top_s1),
      .cpu_data_master_read                                                        (cpu_data_master_read),
      .cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1                       (cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1),
      .cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register        (cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register),
      .cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register             (cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register),
      .cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register              (cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register),
      .cpu_data_master_requests_pb_cpu_to_ddr3_top_s1                              (cpu_data_master_requests_pb_cpu_to_ddr3_top_s1),
      .cpu_data_master_write                                                       (cpu_data_master_write),
      .cpu_data_master_writedata                                                   (cpu_data_master_writedata),
      .cpu_instruction_master_address_to_slave                                     (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1                        (cpu_instruction_master_granted_pb_cpu_to_ddr3_top_s1),
      .cpu_instruction_master_latency_counter                                      (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_pb_cpu_to_ddr3_top_s1              (cpu_instruction_master_qualified_request_pb_cpu_to_ddr3_top_s1),
      .cpu_instruction_master_read                                                 (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1                (cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1),
      .cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register (cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register),
      .cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register      (cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register),
      .cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1                       (cpu_instruction_master_requests_pb_cpu_to_ddr3_top_s1),
      .d1_pb_cpu_to_ddr3_top_s1_end_xfer                                           (d1_pb_cpu_to_ddr3_top_s1_end_xfer),
      .pb_cpu_to_ddr3_top_s1_address                                               (pb_cpu_to_ddr3_top_s1_address),
      .pb_cpu_to_ddr3_top_s1_arbiterlock                                           (pb_cpu_to_ddr3_top_s1_arbiterlock),
      .pb_cpu_to_ddr3_top_s1_arbiterlock2                                          (pb_cpu_to_ddr3_top_s1_arbiterlock2),
      .pb_cpu_to_ddr3_top_s1_burstcount                                            (pb_cpu_to_ddr3_top_s1_burstcount),
      .pb_cpu_to_ddr3_top_s1_byteenable                                            (pb_cpu_to_ddr3_top_s1_byteenable),
      .pb_cpu_to_ddr3_top_s1_chipselect                                            (pb_cpu_to_ddr3_top_s1_chipselect),
      .pb_cpu_to_ddr3_top_s1_debugaccess                                           (pb_cpu_to_ddr3_top_s1_debugaccess),
      .pb_cpu_to_ddr3_top_s1_endofpacket                                           (pb_cpu_to_ddr3_top_s1_endofpacket),
      .pb_cpu_to_ddr3_top_s1_endofpacket_from_sa                                   (pb_cpu_to_ddr3_top_s1_endofpacket_from_sa),
      .pb_cpu_to_ddr3_top_s1_nativeaddress                                         (pb_cpu_to_ddr3_top_s1_nativeaddress),
      .pb_cpu_to_ddr3_top_s1_read                                                  (pb_cpu_to_ddr3_top_s1_read),
      .pb_cpu_to_ddr3_top_s1_readdata                                              (pb_cpu_to_ddr3_top_s1_readdata),
      .pb_cpu_to_ddr3_top_s1_readdata_from_sa                                      (pb_cpu_to_ddr3_top_s1_readdata_from_sa),
      .pb_cpu_to_ddr3_top_s1_readdatavalid                                         (pb_cpu_to_ddr3_top_s1_readdatavalid),
      .pb_cpu_to_ddr3_top_s1_reset_n                                               (pb_cpu_to_ddr3_top_s1_reset_n),
      .pb_cpu_to_ddr3_top_s1_waitrequest                                           (pb_cpu_to_ddr3_top_s1_waitrequest),
      .pb_cpu_to_ddr3_top_s1_waitrequest_from_sa                                   (pb_cpu_to_ddr3_top_s1_waitrequest_from_sa),
      .pb_cpu_to_ddr3_top_s1_write                                                 (pb_cpu_to_ddr3_top_s1_write),
      .pb_cpu_to_ddr3_top_s1_writedata                                             (pb_cpu_to_ddr3_top_s1_writedata),
      .reset_n                                                                     (ddr3_top_phy_clk_out_reset_n)
    );

  pb_cpu_to_ddr3_top_m1_arbitrator the_pb_cpu_to_ddr3_top_m1
    (
      .clk                                                              (ddr3_top_phy_clk_out),
      .d1_ddr3_top_s1_end_xfer                                          (d1_ddr3_top_s1_end_xfer),
      .ddr3_top_s1_readdata_from_sa                                     (ddr3_top_s1_readdata_from_sa),
      .ddr3_top_s1_waitrequest_n_from_sa                                (ddr3_top_s1_waitrequest_n_from_sa),
      .pb_cpu_to_ddr3_top_m1_address                                    (pb_cpu_to_ddr3_top_m1_address),
      .pb_cpu_to_ddr3_top_m1_address_to_slave                           (pb_cpu_to_ddr3_top_m1_address_to_slave),
      .pb_cpu_to_ddr3_top_m1_burstcount                                 (pb_cpu_to_ddr3_top_m1_burstcount),
      .pb_cpu_to_ddr3_top_m1_byteenable                                 (pb_cpu_to_ddr3_top_m1_byteenable),
      .pb_cpu_to_ddr3_top_m1_chipselect                                 (pb_cpu_to_ddr3_top_m1_chipselect),
      .pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1                        (pb_cpu_to_ddr3_top_m1_granted_ddr3_top_s1),
      .pb_cpu_to_ddr3_top_m1_latency_counter                            (pb_cpu_to_ddr3_top_m1_latency_counter),
      .pb_cpu_to_ddr3_top_m1_qualified_request_ddr3_top_s1              (pb_cpu_to_ddr3_top_m1_qualified_request_ddr3_top_s1),
      .pb_cpu_to_ddr3_top_m1_read                                       (pb_cpu_to_ddr3_top_m1_read),
      .pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1                (pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1),
      .pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register (pb_cpu_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register),
      .pb_cpu_to_ddr3_top_m1_readdata                                   (pb_cpu_to_ddr3_top_m1_readdata),
      .pb_cpu_to_ddr3_top_m1_readdatavalid                              (pb_cpu_to_ddr3_top_m1_readdatavalid),
      .pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1                       (pb_cpu_to_ddr3_top_m1_requests_ddr3_top_s1),
      .pb_cpu_to_ddr3_top_m1_waitrequest                                (pb_cpu_to_ddr3_top_m1_waitrequest),
      .pb_cpu_to_ddr3_top_m1_write                                      (pb_cpu_to_ddr3_top_m1_write),
      .pb_cpu_to_ddr3_top_m1_writedata                                  (pb_cpu_to_ddr3_top_m1_writedata),
      .reset_n                                                          (ddr3_top_phy_clk_out_reset_n)
    );

  pb_cpu_to_ddr3_top the_pb_cpu_to_ddr3_top
    (
      .clk              (ddr3_top_phy_clk_out),
      .m1_address       (pb_cpu_to_ddr3_top_m1_address),
      .m1_burstcount    (pb_cpu_to_ddr3_top_m1_burstcount),
      .m1_byteenable    (pb_cpu_to_ddr3_top_m1_byteenable),
      .m1_chipselect    (pb_cpu_to_ddr3_top_m1_chipselect),
      .m1_debugaccess   (pb_cpu_to_ddr3_top_m1_debugaccess),
      .m1_endofpacket   (pb_cpu_to_ddr3_top_m1_endofpacket),
      .m1_read          (pb_cpu_to_ddr3_top_m1_read),
      .m1_readdata      (pb_cpu_to_ddr3_top_m1_readdata),
      .m1_readdatavalid (pb_cpu_to_ddr3_top_m1_readdatavalid),
      .m1_waitrequest   (pb_cpu_to_ddr3_top_m1_waitrequest),
      .m1_write         (pb_cpu_to_ddr3_top_m1_write),
      .m1_writedata     (pb_cpu_to_ddr3_top_m1_writedata),
      .reset_n          (pb_cpu_to_ddr3_top_s1_reset_n),
      .s1_address       (pb_cpu_to_ddr3_top_s1_address),
      .s1_arbiterlock   (pb_cpu_to_ddr3_top_s1_arbiterlock),
      .s1_arbiterlock2  (pb_cpu_to_ddr3_top_s1_arbiterlock2),
      .s1_burstcount    (pb_cpu_to_ddr3_top_s1_burstcount),
      .s1_byteenable    (pb_cpu_to_ddr3_top_s1_byteenable),
      .s1_chipselect    (pb_cpu_to_ddr3_top_s1_chipselect),
      .s1_debugaccess   (pb_cpu_to_ddr3_top_s1_debugaccess),
      .s1_endofpacket   (pb_cpu_to_ddr3_top_s1_endofpacket),
      .s1_nativeaddress (pb_cpu_to_ddr3_top_s1_nativeaddress),
      .s1_read          (pb_cpu_to_ddr3_top_s1_read),
      .s1_readdata      (pb_cpu_to_ddr3_top_s1_readdata),
      .s1_readdatavalid (pb_cpu_to_ddr3_top_s1_readdatavalid),
      .s1_waitrequest   (pb_cpu_to_ddr3_top_s1_waitrequest),
      .s1_write         (pb_cpu_to_ddr3_top_s1_write),
      .s1_writedata     (pb_cpu_to_ddr3_top_s1_writedata)
    );

  pb_cpu_to_fsm_s1_arbitrator the_pb_cpu_to_fsm_s1
    (
      .clk                                                                         (ddr3_top_phy_clk_out),
      .cpu_data_master_address_to_slave                                            (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                  (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                                 (cpu_data_master_debugaccess),
      .cpu_data_master_granted_pb_cpu_to_fsm_s1                                    (cpu_data_master_granted_pb_cpu_to_fsm_s1),
      .cpu_data_master_latency_counter                                             (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_pb_cpu_to_fsm_s1                          (cpu_data_master_qualified_request_pb_cpu_to_fsm_s1),
      .cpu_data_master_read                                                        (cpu_data_master_read),
      .cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register        (cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register),
      .cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1                            (cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1),
      .cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register             (cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register),
      .cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register              (cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register),
      .cpu_data_master_requests_pb_cpu_to_fsm_s1                                   (cpu_data_master_requests_pb_cpu_to_fsm_s1),
      .cpu_data_master_write                                                       (cpu_data_master_write),
      .cpu_data_master_writedata                                                   (cpu_data_master_writedata),
      .cpu_instruction_master_address_to_slave                                     (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_granted_pb_cpu_to_fsm_s1                             (cpu_instruction_master_granted_pb_cpu_to_fsm_s1),
      .cpu_instruction_master_latency_counter                                      (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_pb_cpu_to_fsm_s1                   (cpu_instruction_master_qualified_request_pb_cpu_to_fsm_s1),
      .cpu_instruction_master_read                                                 (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register (cpu_instruction_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register),
      .cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1                     (cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1),
      .cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register      (cpu_instruction_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register),
      .cpu_instruction_master_requests_pb_cpu_to_fsm_s1                            (cpu_instruction_master_requests_pb_cpu_to_fsm_s1),
      .d1_pb_cpu_to_fsm_s1_end_xfer                                                (d1_pb_cpu_to_fsm_s1_end_xfer),
      .pb_cpu_to_fsm_s1_address                                                    (pb_cpu_to_fsm_s1_address),
      .pb_cpu_to_fsm_s1_arbiterlock                                                (pb_cpu_to_fsm_s1_arbiterlock),
      .pb_cpu_to_fsm_s1_arbiterlock2                                               (pb_cpu_to_fsm_s1_arbiterlock2),
      .pb_cpu_to_fsm_s1_burstcount                                                 (pb_cpu_to_fsm_s1_burstcount),
      .pb_cpu_to_fsm_s1_byteenable                                                 (pb_cpu_to_fsm_s1_byteenable),
      .pb_cpu_to_fsm_s1_chipselect                                                 (pb_cpu_to_fsm_s1_chipselect),
      .pb_cpu_to_fsm_s1_debugaccess                                                (pb_cpu_to_fsm_s1_debugaccess),
      .pb_cpu_to_fsm_s1_endofpacket                                                (pb_cpu_to_fsm_s1_endofpacket),
      .pb_cpu_to_fsm_s1_endofpacket_from_sa                                        (pb_cpu_to_fsm_s1_endofpacket_from_sa),
      .pb_cpu_to_fsm_s1_nativeaddress                                              (pb_cpu_to_fsm_s1_nativeaddress),
      .pb_cpu_to_fsm_s1_read                                                       (pb_cpu_to_fsm_s1_read),
      .pb_cpu_to_fsm_s1_readdata                                                   (pb_cpu_to_fsm_s1_readdata),
      .pb_cpu_to_fsm_s1_readdata_from_sa                                           (pb_cpu_to_fsm_s1_readdata_from_sa),
      .pb_cpu_to_fsm_s1_readdatavalid                                              (pb_cpu_to_fsm_s1_readdatavalid),
      .pb_cpu_to_fsm_s1_reset_n                                                    (pb_cpu_to_fsm_s1_reset_n),
      .pb_cpu_to_fsm_s1_waitrequest                                                (pb_cpu_to_fsm_s1_waitrequest),
      .pb_cpu_to_fsm_s1_waitrequest_from_sa                                        (pb_cpu_to_fsm_s1_waitrequest_from_sa),
      .pb_cpu_to_fsm_s1_write                                                      (pb_cpu_to_fsm_s1_write),
      .pb_cpu_to_fsm_s1_writedata                                                  (pb_cpu_to_fsm_s1_writedata),
      .reset_n                                                                     (ddr3_top_phy_clk_out_reset_n)
    );

  pb_cpu_to_fsm_m1_arbitrator the_pb_cpu_to_fsm_m1
    (
      .clk                                               (ddr3_top_phy_clk_out),
      .d1_tb_fsm_avalon_slave_end_xfer                   (d1_tb_fsm_avalon_slave_end_xfer),
      .ext_flash_1_s1_wait_counter_eq_0                  (ext_flash_1_s1_wait_counter_eq_0),
      .ext_flash_s1_wait_counter_eq_0                    (ext_flash_s1_wait_counter_eq_0),
      .incoming_tb_fsm_data_with_Xs_converted_to_0       (incoming_tb_fsm_data_with_Xs_converted_to_0),
      .pb_cpu_to_fsm_m1_address                          (pb_cpu_to_fsm_m1_address),
      .pb_cpu_to_fsm_m1_address_to_slave                 (pb_cpu_to_fsm_m1_address_to_slave),
      .pb_cpu_to_fsm_m1_burstcount                       (pb_cpu_to_fsm_m1_burstcount),
      .pb_cpu_to_fsm_m1_byteenable                       (pb_cpu_to_fsm_m1_byteenable),
      .pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1        (pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1),
      .pb_cpu_to_fsm_m1_byteenable_ext_flash_s1          (pb_cpu_to_fsm_m1_byteenable_ext_flash_s1),
      .pb_cpu_to_fsm_m1_chipselect                       (pb_cpu_to_fsm_m1_chipselect),
      .pb_cpu_to_fsm_m1_dbs_address                      (pb_cpu_to_fsm_m1_dbs_address),
      .pb_cpu_to_fsm_m1_dbs_write_16                     (pb_cpu_to_fsm_m1_dbs_write_16),
      .pb_cpu_to_fsm_m1_granted_ext_flash_1_s1           (pb_cpu_to_fsm_m1_granted_ext_flash_1_s1),
      .pb_cpu_to_fsm_m1_granted_ext_flash_s1             (pb_cpu_to_fsm_m1_granted_ext_flash_s1),
      .pb_cpu_to_fsm_m1_latency_counter                  (pb_cpu_to_fsm_m1_latency_counter),
      .pb_cpu_to_fsm_m1_qualified_request_ext_flash_1_s1 (pb_cpu_to_fsm_m1_qualified_request_ext_flash_1_s1),
      .pb_cpu_to_fsm_m1_qualified_request_ext_flash_s1   (pb_cpu_to_fsm_m1_qualified_request_ext_flash_s1),
      .pb_cpu_to_fsm_m1_read                             (pb_cpu_to_fsm_m1_read),
      .pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1   (pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1),
      .pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1     (pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1),
      .pb_cpu_to_fsm_m1_readdata                         (pb_cpu_to_fsm_m1_readdata),
      .pb_cpu_to_fsm_m1_readdatavalid                    (pb_cpu_to_fsm_m1_readdatavalid),
      .pb_cpu_to_fsm_m1_requests_ext_flash_1_s1          (pb_cpu_to_fsm_m1_requests_ext_flash_1_s1),
      .pb_cpu_to_fsm_m1_requests_ext_flash_s1            (pb_cpu_to_fsm_m1_requests_ext_flash_s1),
      .pb_cpu_to_fsm_m1_waitrequest                      (pb_cpu_to_fsm_m1_waitrequest),
      .pb_cpu_to_fsm_m1_write                            (pb_cpu_to_fsm_m1_write),
      .pb_cpu_to_fsm_m1_writedata                        (pb_cpu_to_fsm_m1_writedata),
      .reset_n                                           (ddr3_top_phy_clk_out_reset_n)
    );

  pb_cpu_to_fsm the_pb_cpu_to_fsm
    (
      .clk              (ddr3_top_phy_clk_out),
      .m1_address       (pb_cpu_to_fsm_m1_address),
      .m1_burstcount    (pb_cpu_to_fsm_m1_burstcount),
      .m1_byteenable    (pb_cpu_to_fsm_m1_byteenable),
      .m1_chipselect    (pb_cpu_to_fsm_m1_chipselect),
      .m1_debugaccess   (pb_cpu_to_fsm_m1_debugaccess),
      .m1_endofpacket   (pb_cpu_to_fsm_m1_endofpacket),
      .m1_read          (pb_cpu_to_fsm_m1_read),
      .m1_readdata      (pb_cpu_to_fsm_m1_readdata),
      .m1_readdatavalid (pb_cpu_to_fsm_m1_readdatavalid),
      .m1_waitrequest   (pb_cpu_to_fsm_m1_waitrequest),
      .m1_write         (pb_cpu_to_fsm_m1_write),
      .m1_writedata     (pb_cpu_to_fsm_m1_writedata),
      .reset_n          (pb_cpu_to_fsm_s1_reset_n),
      .s1_address       (pb_cpu_to_fsm_s1_address),
      .s1_arbiterlock   (pb_cpu_to_fsm_s1_arbiterlock),
      .s1_arbiterlock2  (pb_cpu_to_fsm_s1_arbiterlock2),
      .s1_burstcount    (pb_cpu_to_fsm_s1_burstcount),
      .s1_byteenable    (pb_cpu_to_fsm_s1_byteenable),
      .s1_chipselect    (pb_cpu_to_fsm_s1_chipselect),
      .s1_debugaccess   (pb_cpu_to_fsm_s1_debugaccess),
      .s1_endofpacket   (pb_cpu_to_fsm_s1_endofpacket),
      .s1_nativeaddress (pb_cpu_to_fsm_s1_nativeaddress),
      .s1_read          (pb_cpu_to_fsm_s1_read),
      .s1_readdata      (pb_cpu_to_fsm_s1_readdata),
      .s1_readdatavalid (pb_cpu_to_fsm_s1_readdatavalid),
      .s1_waitrequest   (pb_cpu_to_fsm_s1_waitrequest),
      .s1_write         (pb_cpu_to_fsm_s1_write),
      .s1_writedata     (pb_cpu_to_fsm_s1_writedata)
    );

  pb_cpu_to_io_s1_arbitrator the_pb_cpu_to_io_s1
    (
      .clk                                                                  (ddr3_top_phy_clk_out),
      .cpu_data_master_address_to_slave                                     (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                           (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                          (cpu_data_master_debugaccess),
      .cpu_data_master_granted_pb_cpu_to_io_s1                              (cpu_data_master_granted_pb_cpu_to_io_s1),
      .cpu_data_master_latency_counter                                      (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_pb_cpu_to_io_s1                    (cpu_data_master_qualified_request_pb_cpu_to_io_s1),
      .cpu_data_master_read                                                 (cpu_data_master_read),
      .cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register (cpu_data_master_read_data_valid_pb_cpu_to_ddr3_top_s1_shift_register),
      .cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register      (cpu_data_master_read_data_valid_pb_cpu_to_fsm_s1_shift_register),
      .cpu_data_master_read_data_valid_pb_cpu_to_io_s1                      (cpu_data_master_read_data_valid_pb_cpu_to_io_s1),
      .cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register       (cpu_data_master_read_data_valid_pb_cpu_to_io_s1_shift_register),
      .cpu_data_master_requests_pb_cpu_to_io_s1                             (cpu_data_master_requests_pb_cpu_to_io_s1),
      .cpu_data_master_write                                                (cpu_data_master_write),
      .cpu_data_master_writedata                                            (cpu_data_master_writedata),
      .d1_pb_cpu_to_io_s1_end_xfer                                          (d1_pb_cpu_to_io_s1_end_xfer),
      .pb_cpu_to_io_s1_address                                              (pb_cpu_to_io_s1_address),
      .pb_cpu_to_io_s1_arbiterlock                                          (pb_cpu_to_io_s1_arbiterlock),
      .pb_cpu_to_io_s1_arbiterlock2                                         (pb_cpu_to_io_s1_arbiterlock2),
      .pb_cpu_to_io_s1_burstcount                                           (pb_cpu_to_io_s1_burstcount),
      .pb_cpu_to_io_s1_byteenable                                           (pb_cpu_to_io_s1_byteenable),
      .pb_cpu_to_io_s1_chipselect                                           (pb_cpu_to_io_s1_chipselect),
      .pb_cpu_to_io_s1_debugaccess                                          (pb_cpu_to_io_s1_debugaccess),
      .pb_cpu_to_io_s1_endofpacket                                          (pb_cpu_to_io_s1_endofpacket),
      .pb_cpu_to_io_s1_endofpacket_from_sa                                  (pb_cpu_to_io_s1_endofpacket_from_sa),
      .pb_cpu_to_io_s1_nativeaddress                                        (pb_cpu_to_io_s1_nativeaddress),
      .pb_cpu_to_io_s1_read                                                 (pb_cpu_to_io_s1_read),
      .pb_cpu_to_io_s1_readdata                                             (pb_cpu_to_io_s1_readdata),
      .pb_cpu_to_io_s1_readdata_from_sa                                     (pb_cpu_to_io_s1_readdata_from_sa),
      .pb_cpu_to_io_s1_readdatavalid                                        (pb_cpu_to_io_s1_readdatavalid),
      .pb_cpu_to_io_s1_reset_n                                              (pb_cpu_to_io_s1_reset_n),
      .pb_cpu_to_io_s1_waitrequest                                          (pb_cpu_to_io_s1_waitrequest),
      .pb_cpu_to_io_s1_waitrequest_from_sa                                  (pb_cpu_to_io_s1_waitrequest_from_sa),
      .pb_cpu_to_io_s1_write                                                (pb_cpu_to_io_s1_write),
      .pb_cpu_to_io_s1_writedata                                            (pb_cpu_to_io_s1_writedata),
      .reset_n                                                              (ddr3_top_phy_clk_out_reset_n)
    );

  pb_cpu_to_io_m1_arbitrator the_pb_cpu_to_io_m1
    (
      .button_pio_s1_readdata_from_sa                                (button_pio_s1_readdata_from_sa),
      .clk                                                           (ddr3_top_phy_clk_out),
      .d1_button_pio_s1_end_xfer                                     (d1_button_pio_s1_end_xfer),
      .d1_descriptor_memory_s1_end_xfer                              (d1_descriptor_memory_s1_end_xfer),
      .d1_dipsw_pio_s1_end_xfer                                      (d1_dipsw_pio_s1_end_xfer),
      .d1_jtag_uart_avalon_jtag_slave_end_xfer                       (d1_jtag_uart_avalon_jtag_slave_end_xfer),
      .d1_led_pio_s1_end_xfer                                        (d1_led_pio_s1_end_xfer),
      .d1_sgdma_rx_csr_end_xfer                                      (d1_sgdma_rx_csr_end_xfer),
      .d1_sgdma_tx_csr_end_xfer                                      (d1_sgdma_tx_csr_end_xfer),
      .d1_sysid_control_slave_end_xfer                               (d1_sysid_control_slave_end_xfer),
      .d1_timer_1ms_s1_end_xfer                                      (d1_timer_1ms_s1_end_xfer),
      .d1_tse_mac_control_port_end_xfer                              (d1_tse_mac_control_port_end_xfer),
      .d1_uart_s1_end_xfer                                           (d1_uart_s1_end_xfer),
      .descriptor_memory_s1_readdata_from_sa                         (descriptor_memory_s1_readdata_from_sa),
      .dipsw_pio_s1_readdata_from_sa                                 (dipsw_pio_s1_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_readdata_from_sa                  (jtag_uart_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_waitrequest_from_sa               (jtag_uart_avalon_jtag_slave_waitrequest_from_sa),
      .led_pio_s1_readdata_from_sa                                   (led_pio_s1_readdata_from_sa),
      .pb_cpu_to_io_m1_address                                       (pb_cpu_to_io_m1_address),
      .pb_cpu_to_io_m1_address_to_slave                              (pb_cpu_to_io_m1_address_to_slave),
      .pb_cpu_to_io_m1_burstcount                                    (pb_cpu_to_io_m1_burstcount),
      .pb_cpu_to_io_m1_byteenable                                    (pb_cpu_to_io_m1_byteenable),
      .pb_cpu_to_io_m1_chipselect                                    (pb_cpu_to_io_m1_chipselect),
      .pb_cpu_to_io_m1_granted_button_pio_s1                         (pb_cpu_to_io_m1_granted_button_pio_s1),
      .pb_cpu_to_io_m1_granted_descriptor_memory_s1                  (pb_cpu_to_io_m1_granted_descriptor_memory_s1),
      .pb_cpu_to_io_m1_granted_dipsw_pio_s1                          (pb_cpu_to_io_m1_granted_dipsw_pio_s1),
      .pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave           (pb_cpu_to_io_m1_granted_jtag_uart_avalon_jtag_slave),
      .pb_cpu_to_io_m1_granted_led_pio_s1                            (pb_cpu_to_io_m1_granted_led_pio_s1),
      .pb_cpu_to_io_m1_granted_sgdma_rx_csr                          (pb_cpu_to_io_m1_granted_sgdma_rx_csr),
      .pb_cpu_to_io_m1_granted_sgdma_tx_csr                          (pb_cpu_to_io_m1_granted_sgdma_tx_csr),
      .pb_cpu_to_io_m1_granted_sysid_control_slave                   (pb_cpu_to_io_m1_granted_sysid_control_slave),
      .pb_cpu_to_io_m1_granted_timer_1ms_s1                          (pb_cpu_to_io_m1_granted_timer_1ms_s1),
      .pb_cpu_to_io_m1_granted_tse_mac_control_port                  (pb_cpu_to_io_m1_granted_tse_mac_control_port),
      .pb_cpu_to_io_m1_granted_uart_s1                               (pb_cpu_to_io_m1_granted_uart_s1),
      .pb_cpu_to_io_m1_latency_counter                               (pb_cpu_to_io_m1_latency_counter),
      .pb_cpu_to_io_m1_qualified_request_button_pio_s1               (pb_cpu_to_io_m1_qualified_request_button_pio_s1),
      .pb_cpu_to_io_m1_qualified_request_descriptor_memory_s1        (pb_cpu_to_io_m1_qualified_request_descriptor_memory_s1),
      .pb_cpu_to_io_m1_qualified_request_dipsw_pio_s1                (pb_cpu_to_io_m1_qualified_request_dipsw_pio_s1),
      .pb_cpu_to_io_m1_qualified_request_jtag_uart_avalon_jtag_slave (pb_cpu_to_io_m1_qualified_request_jtag_uart_avalon_jtag_slave),
      .pb_cpu_to_io_m1_qualified_request_led_pio_s1                  (pb_cpu_to_io_m1_qualified_request_led_pio_s1),
      .pb_cpu_to_io_m1_qualified_request_sgdma_rx_csr                (pb_cpu_to_io_m1_qualified_request_sgdma_rx_csr),
      .pb_cpu_to_io_m1_qualified_request_sgdma_tx_csr                (pb_cpu_to_io_m1_qualified_request_sgdma_tx_csr),
      .pb_cpu_to_io_m1_qualified_request_sysid_control_slave         (pb_cpu_to_io_m1_qualified_request_sysid_control_slave),
      .pb_cpu_to_io_m1_qualified_request_timer_1ms_s1                (pb_cpu_to_io_m1_qualified_request_timer_1ms_s1),
      .pb_cpu_to_io_m1_qualified_request_tse_mac_control_port        (pb_cpu_to_io_m1_qualified_request_tse_mac_control_port),
      .pb_cpu_to_io_m1_qualified_request_uart_s1                     (pb_cpu_to_io_m1_qualified_request_uart_s1),
      .pb_cpu_to_io_m1_read                                          (pb_cpu_to_io_m1_read),
      .pb_cpu_to_io_m1_read_data_valid_button_pio_s1                 (pb_cpu_to_io_m1_read_data_valid_button_pio_s1),
      .pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1          (pb_cpu_to_io_m1_read_data_valid_descriptor_memory_s1),
      .pb_cpu_to_io_m1_read_data_valid_dipsw_pio_s1                  (pb_cpu_to_io_m1_read_data_valid_dipsw_pio_s1),
      .pb_cpu_to_io_m1_read_data_valid_jtag_uart_avalon_jtag_slave   (pb_cpu_to_io_m1_read_data_valid_jtag_uart_avalon_jtag_slave),
      .pb_cpu_to_io_m1_read_data_valid_led_pio_s1                    (pb_cpu_to_io_m1_read_data_valid_led_pio_s1),
      .pb_cpu_to_io_m1_read_data_valid_sgdma_rx_csr                  (pb_cpu_to_io_m1_read_data_valid_sgdma_rx_csr),
      .pb_cpu_to_io_m1_read_data_valid_sgdma_tx_csr                  (pb_cpu_to_io_m1_read_data_valid_sgdma_tx_csr),
      .pb_cpu_to_io_m1_read_data_valid_sysid_control_slave           (pb_cpu_to_io_m1_read_data_valid_sysid_control_slave),
      .pb_cpu_to_io_m1_read_data_valid_timer_1ms_s1                  (pb_cpu_to_io_m1_read_data_valid_timer_1ms_s1),
      .pb_cpu_to_io_m1_read_data_valid_tse_mac_control_port          (pb_cpu_to_io_m1_read_data_valid_tse_mac_control_port),
      .pb_cpu_to_io_m1_read_data_valid_uart_s1                       (pb_cpu_to_io_m1_read_data_valid_uart_s1),
      .pb_cpu_to_io_m1_readdata                                      (pb_cpu_to_io_m1_readdata),
      .pb_cpu_to_io_m1_readdatavalid                                 (pb_cpu_to_io_m1_readdatavalid),
      .pb_cpu_to_io_m1_requests_button_pio_s1                        (pb_cpu_to_io_m1_requests_button_pio_s1),
      .pb_cpu_to_io_m1_requests_descriptor_memory_s1                 (pb_cpu_to_io_m1_requests_descriptor_memory_s1),
      .pb_cpu_to_io_m1_requests_dipsw_pio_s1                         (pb_cpu_to_io_m1_requests_dipsw_pio_s1),
      .pb_cpu_to_io_m1_requests_jtag_uart_avalon_jtag_slave          (pb_cpu_to_io_m1_requests_jtag_uart_avalon_jtag_slave),
      .pb_cpu_to_io_m1_requests_led_pio_s1                           (pb_cpu_to_io_m1_requests_led_pio_s1),
      .pb_cpu_to_io_m1_requests_sgdma_rx_csr                         (pb_cpu_to_io_m1_requests_sgdma_rx_csr),
      .pb_cpu_to_io_m1_requests_sgdma_tx_csr                         (pb_cpu_to_io_m1_requests_sgdma_tx_csr),
      .pb_cpu_to_io_m1_requests_sysid_control_slave                  (pb_cpu_to_io_m1_requests_sysid_control_slave),
      .pb_cpu_to_io_m1_requests_timer_1ms_s1                         (pb_cpu_to_io_m1_requests_timer_1ms_s1),
      .pb_cpu_to_io_m1_requests_tse_mac_control_port                 (pb_cpu_to_io_m1_requests_tse_mac_control_port),
      .pb_cpu_to_io_m1_requests_uart_s1                              (pb_cpu_to_io_m1_requests_uart_s1),
      .pb_cpu_to_io_m1_waitrequest                                   (pb_cpu_to_io_m1_waitrequest),
      .pb_cpu_to_io_m1_write                                         (pb_cpu_to_io_m1_write),
      .pb_cpu_to_io_m1_writedata                                     (pb_cpu_to_io_m1_writedata),
      .reset_n                                                       (ddr3_top_phy_clk_out_reset_n),
      .sgdma_rx_csr_readdata_from_sa                                 (sgdma_rx_csr_readdata_from_sa),
      .sgdma_tx_csr_readdata_from_sa                                 (sgdma_tx_csr_readdata_from_sa),
      .sysid_control_slave_readdata_from_sa                          (sysid_control_slave_readdata_from_sa),
      .timer_1ms_s1_readdata_from_sa                                 (timer_1ms_s1_readdata_from_sa),
      .tse_mac_control_port_readdata_from_sa                         (tse_mac_control_port_readdata_from_sa),
      .tse_mac_control_port_waitrequest_from_sa                      (tse_mac_control_port_waitrequest_from_sa),
      .uart_s1_readdata_from_sa                                      (uart_s1_readdata_from_sa)
    );

  pb_cpu_to_io the_pb_cpu_to_io
    (
      .clk              (ddr3_top_phy_clk_out),
      .m1_address       (pb_cpu_to_io_m1_address),
      .m1_burstcount    (pb_cpu_to_io_m1_burstcount),
      .m1_byteenable    (pb_cpu_to_io_m1_byteenable),
      .m1_chipselect    (pb_cpu_to_io_m1_chipselect),
      .m1_debugaccess   (pb_cpu_to_io_m1_debugaccess),
      .m1_endofpacket   (pb_cpu_to_io_m1_endofpacket),
      .m1_read          (pb_cpu_to_io_m1_read),
      .m1_readdata      (pb_cpu_to_io_m1_readdata),
      .m1_readdatavalid (pb_cpu_to_io_m1_readdatavalid),
      .m1_waitrequest   (pb_cpu_to_io_m1_waitrequest),
      .m1_write         (pb_cpu_to_io_m1_write),
      .m1_writedata     (pb_cpu_to_io_m1_writedata),
      .reset_n          (pb_cpu_to_io_s1_reset_n),
      .s1_address       (pb_cpu_to_io_s1_address),
      .s1_arbiterlock   (pb_cpu_to_io_s1_arbiterlock),
      .s1_arbiterlock2  (pb_cpu_to_io_s1_arbiterlock2),
      .s1_burstcount    (pb_cpu_to_io_s1_burstcount),
      .s1_byteenable    (pb_cpu_to_io_s1_byteenable),
      .s1_chipselect    (pb_cpu_to_io_s1_chipselect),
      .s1_debugaccess   (pb_cpu_to_io_s1_debugaccess),
      .s1_endofpacket   (pb_cpu_to_io_s1_endofpacket),
      .s1_nativeaddress (pb_cpu_to_io_s1_nativeaddress),
      .s1_read          (pb_cpu_to_io_s1_read),
      .s1_readdata      (pb_cpu_to_io_s1_readdata),
      .s1_readdatavalid (pb_cpu_to_io_s1_readdatavalid),
      .s1_waitrequest   (pb_cpu_to_io_s1_waitrequest),
      .s1_write         (pb_cpu_to_io_s1_write),
      .s1_writedata     (pb_cpu_to_io_s1_writedata)
    );

  pb_dma_to_ddr3_top_s1_arbitrator the_pb_dma_to_ddr3_top_s1
    (
      .clk                                                                  (ddr3_top_phy_clk_out),
      .d1_pb_dma_to_ddr3_top_s1_end_xfer                                    (d1_pb_dma_to_ddr3_top_s1_end_xfer),
      .pb_dma_to_ddr3_top_s1_address                                        (pb_dma_to_ddr3_top_s1_address),
      .pb_dma_to_ddr3_top_s1_arbiterlock                                    (pb_dma_to_ddr3_top_s1_arbiterlock),
      .pb_dma_to_ddr3_top_s1_arbiterlock2                                   (pb_dma_to_ddr3_top_s1_arbiterlock2),
      .pb_dma_to_ddr3_top_s1_burstcount                                     (pb_dma_to_ddr3_top_s1_burstcount),
      .pb_dma_to_ddr3_top_s1_byteenable                                     (pb_dma_to_ddr3_top_s1_byteenable),
      .pb_dma_to_ddr3_top_s1_chipselect                                     (pb_dma_to_ddr3_top_s1_chipselect),
      .pb_dma_to_ddr3_top_s1_debugaccess                                    (pb_dma_to_ddr3_top_s1_debugaccess),
      .pb_dma_to_ddr3_top_s1_endofpacket                                    (pb_dma_to_ddr3_top_s1_endofpacket),
      .pb_dma_to_ddr3_top_s1_endofpacket_from_sa                            (pb_dma_to_ddr3_top_s1_endofpacket_from_sa),
      .pb_dma_to_ddr3_top_s1_nativeaddress                                  (pb_dma_to_ddr3_top_s1_nativeaddress),
      .pb_dma_to_ddr3_top_s1_read                                           (pb_dma_to_ddr3_top_s1_read),
      .pb_dma_to_ddr3_top_s1_readdata                                       (pb_dma_to_ddr3_top_s1_readdata),
      .pb_dma_to_ddr3_top_s1_readdata_from_sa                               (pb_dma_to_ddr3_top_s1_readdata_from_sa),
      .pb_dma_to_ddr3_top_s1_readdatavalid                                  (pb_dma_to_ddr3_top_s1_readdatavalid),
      .pb_dma_to_ddr3_top_s1_reset_n                                        (pb_dma_to_ddr3_top_s1_reset_n),
      .pb_dma_to_ddr3_top_s1_waitrequest                                    (pb_dma_to_ddr3_top_s1_waitrequest),
      .pb_dma_to_ddr3_top_s1_waitrequest_from_sa                            (pb_dma_to_ddr3_top_s1_waitrequest_from_sa),
      .pb_dma_to_ddr3_top_s1_write                                          (pb_dma_to_ddr3_top_s1_write),
      .pb_dma_to_ddr3_top_s1_writedata                                      (pb_dma_to_ddr3_top_s1_writedata),
      .reset_n                                                              (ddr3_top_phy_clk_out_reset_n),
      .sgdma_rx_m_write_address_to_slave                                    (sgdma_rx_m_write_address_to_slave),
      .sgdma_rx_m_write_byteenable                                          (sgdma_rx_m_write_byteenable),
      .sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1                       (sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1),
      .sgdma_rx_m_write_qualified_request_pb_dma_to_ddr3_top_s1             (sgdma_rx_m_write_qualified_request_pb_dma_to_ddr3_top_s1),
      .sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1                      (sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1),
      .sgdma_rx_m_write_write                                               (sgdma_rx_m_write_write),
      .sgdma_rx_m_write_writedata                                           (sgdma_rx_m_write_writedata),
      .sgdma_tx_m_read_address_to_slave                                     (sgdma_tx_m_read_address_to_slave),
      .sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1                        (sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1),
      .sgdma_tx_m_read_latency_counter                                      (sgdma_tx_m_read_latency_counter),
      .sgdma_tx_m_read_qualified_request_pb_dma_to_ddr3_top_s1              (sgdma_tx_m_read_qualified_request_pb_dma_to_ddr3_top_s1),
      .sgdma_tx_m_read_read                                                 (sgdma_tx_m_read_read),
      .sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1                (sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1),
      .sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1_shift_register (sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1_shift_register),
      .sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1                       (sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1)
    );

  pb_dma_to_ddr3_top_m1_arbitrator the_pb_dma_to_ddr3_top_m1
    (
      .clk                                                              (ddr3_top_phy_clk_out),
      .d1_ddr3_top_s1_end_xfer                                          (d1_ddr3_top_s1_end_xfer),
      .ddr3_top_s1_readdata_from_sa                                     (ddr3_top_s1_readdata_from_sa),
      .ddr3_top_s1_waitrequest_n_from_sa                                (ddr3_top_s1_waitrequest_n_from_sa),
      .pb_dma_to_ddr3_top_m1_address                                    (pb_dma_to_ddr3_top_m1_address),
      .pb_dma_to_ddr3_top_m1_address_to_slave                           (pb_dma_to_ddr3_top_m1_address_to_slave),
      .pb_dma_to_ddr3_top_m1_burstcount                                 (pb_dma_to_ddr3_top_m1_burstcount),
      .pb_dma_to_ddr3_top_m1_byteenable                                 (pb_dma_to_ddr3_top_m1_byteenable),
      .pb_dma_to_ddr3_top_m1_chipselect                                 (pb_dma_to_ddr3_top_m1_chipselect),
      .pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1                        (pb_dma_to_ddr3_top_m1_granted_ddr3_top_s1),
      .pb_dma_to_ddr3_top_m1_latency_counter                            (pb_dma_to_ddr3_top_m1_latency_counter),
      .pb_dma_to_ddr3_top_m1_qualified_request_ddr3_top_s1              (pb_dma_to_ddr3_top_m1_qualified_request_ddr3_top_s1),
      .pb_dma_to_ddr3_top_m1_read                                       (pb_dma_to_ddr3_top_m1_read),
      .pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1                (pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1),
      .pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register (pb_dma_to_ddr3_top_m1_read_data_valid_ddr3_top_s1_shift_register),
      .pb_dma_to_ddr3_top_m1_readdata                                   (pb_dma_to_ddr3_top_m1_readdata),
      .pb_dma_to_ddr3_top_m1_readdatavalid                              (pb_dma_to_ddr3_top_m1_readdatavalid),
      .pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1                       (pb_dma_to_ddr3_top_m1_requests_ddr3_top_s1),
      .pb_dma_to_ddr3_top_m1_waitrequest                                (pb_dma_to_ddr3_top_m1_waitrequest),
      .pb_dma_to_ddr3_top_m1_write                                      (pb_dma_to_ddr3_top_m1_write),
      .pb_dma_to_ddr3_top_m1_writedata                                  (pb_dma_to_ddr3_top_m1_writedata),
      .reset_n                                                          (ddr3_top_phy_clk_out_reset_n)
    );

  pb_dma_to_ddr3_top the_pb_dma_to_ddr3_top
    (
      .clk              (ddr3_top_phy_clk_out),
      .m1_address       (pb_dma_to_ddr3_top_m1_address),
      .m1_burstcount    (pb_dma_to_ddr3_top_m1_burstcount),
      .m1_byteenable    (pb_dma_to_ddr3_top_m1_byteenable),
      .m1_chipselect    (pb_dma_to_ddr3_top_m1_chipselect),
      .m1_debugaccess   (pb_dma_to_ddr3_top_m1_debugaccess),
      .m1_endofpacket   (pb_dma_to_ddr3_top_m1_endofpacket),
      .m1_read          (pb_dma_to_ddr3_top_m1_read),
      .m1_readdata      (pb_dma_to_ddr3_top_m1_readdata),
      .m1_readdatavalid (pb_dma_to_ddr3_top_m1_readdatavalid),
      .m1_waitrequest   (pb_dma_to_ddr3_top_m1_waitrequest),
      .m1_write         (pb_dma_to_ddr3_top_m1_write),
      .m1_writedata     (pb_dma_to_ddr3_top_m1_writedata),
      .reset_n          (pb_dma_to_ddr3_top_s1_reset_n),
      .s1_address       (pb_dma_to_ddr3_top_s1_address),
      .s1_arbiterlock   (pb_dma_to_ddr3_top_s1_arbiterlock),
      .s1_arbiterlock2  (pb_dma_to_ddr3_top_s1_arbiterlock2),
      .s1_burstcount    (pb_dma_to_ddr3_top_s1_burstcount),
      .s1_byteenable    (pb_dma_to_ddr3_top_s1_byteenable),
      .s1_chipselect    (pb_dma_to_ddr3_top_s1_chipselect),
      .s1_debugaccess   (pb_dma_to_ddr3_top_s1_debugaccess),
      .s1_endofpacket   (pb_dma_to_ddr3_top_s1_endofpacket),
      .s1_nativeaddress (pb_dma_to_ddr3_top_s1_nativeaddress),
      .s1_read          (pb_dma_to_ddr3_top_s1_read),
      .s1_readdata      (pb_dma_to_ddr3_top_s1_readdata),
      .s1_readdatavalid (pb_dma_to_ddr3_top_s1_readdatavalid),
      .s1_waitrequest   (pb_dma_to_ddr3_top_s1_waitrequest),
      .s1_write         (pb_dma_to_ddr3_top_s1_write),
      .s1_writedata     (pb_dma_to_ddr3_top_s1_writedata)
    );

  pb_dma_to_descriptor_memory_s1_arbitrator the_pb_dma_to_descriptor_memory_s1
    (
      .clk                                                                                    (ddr3_top_phy_clk_out),
      .d1_pb_dma_to_descriptor_memory_s1_end_xfer                                             (d1_pb_dma_to_descriptor_memory_s1_end_xfer),
      .pb_dma_to_descriptor_memory_s1_address                                                 (pb_dma_to_descriptor_memory_s1_address),
      .pb_dma_to_descriptor_memory_s1_arbiterlock                                             (pb_dma_to_descriptor_memory_s1_arbiterlock),
      .pb_dma_to_descriptor_memory_s1_arbiterlock2                                            (pb_dma_to_descriptor_memory_s1_arbiterlock2),
      .pb_dma_to_descriptor_memory_s1_burstcount                                              (pb_dma_to_descriptor_memory_s1_burstcount),
      .pb_dma_to_descriptor_memory_s1_byteenable                                              (pb_dma_to_descriptor_memory_s1_byteenable),
      .pb_dma_to_descriptor_memory_s1_chipselect                                              (pb_dma_to_descriptor_memory_s1_chipselect),
      .pb_dma_to_descriptor_memory_s1_debugaccess                                             (pb_dma_to_descriptor_memory_s1_debugaccess),
      .pb_dma_to_descriptor_memory_s1_endofpacket                                             (pb_dma_to_descriptor_memory_s1_endofpacket),
      .pb_dma_to_descriptor_memory_s1_endofpacket_from_sa                                     (pb_dma_to_descriptor_memory_s1_endofpacket_from_sa),
      .pb_dma_to_descriptor_memory_s1_nativeaddress                                           (pb_dma_to_descriptor_memory_s1_nativeaddress),
      .pb_dma_to_descriptor_memory_s1_read                                                    (pb_dma_to_descriptor_memory_s1_read),
      .pb_dma_to_descriptor_memory_s1_readdata                                                (pb_dma_to_descriptor_memory_s1_readdata),
      .pb_dma_to_descriptor_memory_s1_readdata_from_sa                                        (pb_dma_to_descriptor_memory_s1_readdata_from_sa),
      .pb_dma_to_descriptor_memory_s1_readdatavalid                                           (pb_dma_to_descriptor_memory_s1_readdatavalid),
      .pb_dma_to_descriptor_memory_s1_reset_n                                                 (pb_dma_to_descriptor_memory_s1_reset_n),
      .pb_dma_to_descriptor_memory_s1_waitrequest                                             (pb_dma_to_descriptor_memory_s1_waitrequest),
      .pb_dma_to_descriptor_memory_s1_waitrequest_from_sa                                     (pb_dma_to_descriptor_memory_s1_waitrequest_from_sa),
      .pb_dma_to_descriptor_memory_s1_write                                                   (pb_dma_to_descriptor_memory_s1_write),
      .pb_dma_to_descriptor_memory_s1_writedata                                               (pb_dma_to_descriptor_memory_s1_writedata),
      .reset_n                                                                                (ddr3_top_phy_clk_out_reset_n),
      .sgdma_rx_descriptor_read_address_to_slave                                              (sgdma_rx_descriptor_read_address_to_slave),
      .sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1                        (sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_latency_counter                                               (sgdma_rx_descriptor_read_latency_counter),
      .sgdma_rx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1              (sgdma_rx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_read                                                          (sgdma_rx_descriptor_read_read),
      .sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1                (sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register (sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register),
      .sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1                       (sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_address_to_slave                                             (sgdma_rx_descriptor_write_address_to_slave),
      .sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1                       (sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1             (sgdma_rx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1                      (sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_write                                                        (sgdma_rx_descriptor_write_write),
      .sgdma_rx_descriptor_write_writedata                                                    (sgdma_rx_descriptor_write_writedata),
      .sgdma_tx_descriptor_read_address_to_slave                                              (sgdma_tx_descriptor_read_address_to_slave),
      .sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1                        (sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_latency_counter                                               (sgdma_tx_descriptor_read_latency_counter),
      .sgdma_tx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1              (sgdma_tx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_read                                                          (sgdma_tx_descriptor_read_read),
      .sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1                (sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register (sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register),
      .sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1                       (sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_address_to_slave                                             (sgdma_tx_descriptor_write_address_to_slave),
      .sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1                       (sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1             (sgdma_tx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1                      (sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_write                                                        (sgdma_tx_descriptor_write_write),
      .sgdma_tx_descriptor_write_writedata                                                    (sgdma_tx_descriptor_write_writedata)
    );

  pb_dma_to_descriptor_memory_m1_arbitrator the_pb_dma_to_descriptor_memory_m1
    (
      .clk                                                                   (ddr3_top_phy_clk_out),
      .d1_descriptor_memory_s1_end_xfer                                      (d1_descriptor_memory_s1_end_xfer),
      .descriptor_memory_s1_readdata_from_sa                                 (descriptor_memory_s1_readdata_from_sa),
      .pb_dma_to_descriptor_memory_m1_address                                (pb_dma_to_descriptor_memory_m1_address),
      .pb_dma_to_descriptor_memory_m1_address_to_slave                       (pb_dma_to_descriptor_memory_m1_address_to_slave),
      .pb_dma_to_descriptor_memory_m1_burstcount                             (pb_dma_to_descriptor_memory_m1_burstcount),
      .pb_dma_to_descriptor_memory_m1_byteenable                             (pb_dma_to_descriptor_memory_m1_byteenable),
      .pb_dma_to_descriptor_memory_m1_chipselect                             (pb_dma_to_descriptor_memory_m1_chipselect),
      .pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1           (pb_dma_to_descriptor_memory_m1_granted_descriptor_memory_s1),
      .pb_dma_to_descriptor_memory_m1_latency_counter                        (pb_dma_to_descriptor_memory_m1_latency_counter),
      .pb_dma_to_descriptor_memory_m1_qualified_request_descriptor_memory_s1 (pb_dma_to_descriptor_memory_m1_qualified_request_descriptor_memory_s1),
      .pb_dma_to_descriptor_memory_m1_read                                   (pb_dma_to_descriptor_memory_m1_read),
      .pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1   (pb_dma_to_descriptor_memory_m1_read_data_valid_descriptor_memory_s1),
      .pb_dma_to_descriptor_memory_m1_readdata                               (pb_dma_to_descriptor_memory_m1_readdata),
      .pb_dma_to_descriptor_memory_m1_readdatavalid                          (pb_dma_to_descriptor_memory_m1_readdatavalid),
      .pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1          (pb_dma_to_descriptor_memory_m1_requests_descriptor_memory_s1),
      .pb_dma_to_descriptor_memory_m1_waitrequest                            (pb_dma_to_descriptor_memory_m1_waitrequest),
      .pb_dma_to_descriptor_memory_m1_write                                  (pb_dma_to_descriptor_memory_m1_write),
      .pb_dma_to_descriptor_memory_m1_writedata                              (pb_dma_to_descriptor_memory_m1_writedata),
      .reset_n                                                               (ddr3_top_phy_clk_out_reset_n)
    );

  pb_dma_to_descriptor_memory the_pb_dma_to_descriptor_memory
    (
      .clk              (ddr3_top_phy_clk_out),
      .m1_address       (pb_dma_to_descriptor_memory_m1_address),
      .m1_burstcount    (pb_dma_to_descriptor_memory_m1_burstcount),
      .m1_byteenable    (pb_dma_to_descriptor_memory_m1_byteenable),
      .m1_chipselect    (pb_dma_to_descriptor_memory_m1_chipselect),
      .m1_debugaccess   (pb_dma_to_descriptor_memory_m1_debugaccess),
      .m1_endofpacket   (pb_dma_to_descriptor_memory_m1_endofpacket),
      .m1_read          (pb_dma_to_descriptor_memory_m1_read),
      .m1_readdata      (pb_dma_to_descriptor_memory_m1_readdata),
      .m1_readdatavalid (pb_dma_to_descriptor_memory_m1_readdatavalid),
      .m1_waitrequest   (pb_dma_to_descriptor_memory_m1_waitrequest),
      .m1_write         (pb_dma_to_descriptor_memory_m1_write),
      .m1_writedata     (pb_dma_to_descriptor_memory_m1_writedata),
      .reset_n          (pb_dma_to_descriptor_memory_s1_reset_n),
      .s1_address       (pb_dma_to_descriptor_memory_s1_address),
      .s1_arbiterlock   (pb_dma_to_descriptor_memory_s1_arbiterlock),
      .s1_arbiterlock2  (pb_dma_to_descriptor_memory_s1_arbiterlock2),
      .s1_burstcount    (pb_dma_to_descriptor_memory_s1_burstcount),
      .s1_byteenable    (pb_dma_to_descriptor_memory_s1_byteenable),
      .s1_chipselect    (pb_dma_to_descriptor_memory_s1_chipselect),
      .s1_debugaccess   (pb_dma_to_descriptor_memory_s1_debugaccess),
      .s1_endofpacket   (pb_dma_to_descriptor_memory_s1_endofpacket),
      .s1_nativeaddress (pb_dma_to_descriptor_memory_s1_nativeaddress),
      .s1_read          (pb_dma_to_descriptor_memory_s1_read),
      .s1_readdata      (pb_dma_to_descriptor_memory_s1_readdata),
      .s1_readdatavalid (pb_dma_to_descriptor_memory_s1_readdatavalid),
      .s1_waitrequest   (pb_dma_to_descriptor_memory_s1_waitrequest),
      .s1_write         (pb_dma_to_descriptor_memory_s1_write),
      .s1_writedata     (pb_dma_to_descriptor_memory_s1_writedata)
    );

  sgdma_rx_csr_arbitrator the_sgdma_rx_csr
    (
      .clk                                            (ddr3_top_phy_clk_out),
      .d1_sgdma_rx_csr_end_xfer                       (d1_sgdma_rx_csr_end_xfer),
      .pb_cpu_to_io_m1_address_to_slave               (pb_cpu_to_io_m1_address_to_slave),
      .pb_cpu_to_io_m1_burstcount                     (pb_cpu_to_io_m1_burstcount),
      .pb_cpu_to_io_m1_chipselect                     (pb_cpu_to_io_m1_chipselect),
      .pb_cpu_to_io_m1_granted_sgdma_rx_csr           (pb_cpu_to_io_m1_granted_sgdma_rx_csr),
      .pb_cpu_to_io_m1_latency_counter                (pb_cpu_to_io_m1_latency_counter),
      .pb_cpu_to_io_m1_qualified_request_sgdma_rx_csr (pb_cpu_to_io_m1_qualified_request_sgdma_rx_csr),
      .pb_cpu_to_io_m1_read                           (pb_cpu_to_io_m1_read),
      .pb_cpu_to_io_m1_read_data_valid_sgdma_rx_csr   (pb_cpu_to_io_m1_read_data_valid_sgdma_rx_csr),
      .pb_cpu_to_io_m1_requests_sgdma_rx_csr          (pb_cpu_to_io_m1_requests_sgdma_rx_csr),
      .pb_cpu_to_io_m1_write                          (pb_cpu_to_io_m1_write),
      .pb_cpu_to_io_m1_writedata                      (pb_cpu_to_io_m1_writedata),
      .reset_n                                        (ddr3_top_phy_clk_out_reset_n),
      .sgdma_rx_csr_address                           (sgdma_rx_csr_address),
      .sgdma_rx_csr_chipselect                        (sgdma_rx_csr_chipselect),
      .sgdma_rx_csr_irq                               (sgdma_rx_csr_irq),
      .sgdma_rx_csr_irq_from_sa                       (sgdma_rx_csr_irq_from_sa),
      .sgdma_rx_csr_read                              (sgdma_rx_csr_read),
      .sgdma_rx_csr_readdata                          (sgdma_rx_csr_readdata),
      .sgdma_rx_csr_readdata_from_sa                  (sgdma_rx_csr_readdata_from_sa),
      .sgdma_rx_csr_reset_n                           (sgdma_rx_csr_reset_n),
      .sgdma_rx_csr_write                             (sgdma_rx_csr_write),
      .sgdma_rx_csr_writedata                         (sgdma_rx_csr_writedata)
    );

  sgdma_rx_in_arbitrator the_sgdma_rx_in
    (
      .clk                           (ddr3_top_phy_clk_out),
      .reset_n                       (ddr3_top_phy_clk_out_reset_n),
      .sgdma_rx_in_data              (sgdma_rx_in_data),
      .sgdma_rx_in_empty             (sgdma_rx_in_empty),
      .sgdma_rx_in_endofpacket       (sgdma_rx_in_endofpacket),
      .sgdma_rx_in_error             (sgdma_rx_in_error),
      .sgdma_rx_in_ready             (sgdma_rx_in_ready),
      .sgdma_rx_in_ready_from_sa     (sgdma_rx_in_ready_from_sa),
      .sgdma_rx_in_startofpacket     (sgdma_rx_in_startofpacket),
      .sgdma_rx_in_valid             (sgdma_rx_in_valid),
      .tse_mac_receive_data          (tse_mac_receive_data),
      .tse_mac_receive_empty         (tse_mac_receive_empty),
      .tse_mac_receive_endofpacket   (tse_mac_receive_endofpacket),
      .tse_mac_receive_error         (tse_mac_receive_error),
      .tse_mac_receive_startofpacket (tse_mac_receive_startofpacket),
      .tse_mac_receive_valid         (tse_mac_receive_valid)
    );

  sgdma_rx_descriptor_read_arbitrator the_sgdma_rx_descriptor_read
    (
      .clk                                                                                    (ddr3_top_phy_clk_out),
      .d1_pb_dma_to_descriptor_memory_s1_end_xfer                                             (d1_pb_dma_to_descriptor_memory_s1_end_xfer),
      .pb_dma_to_descriptor_memory_s1_readdata_from_sa                                        (pb_dma_to_descriptor_memory_s1_readdata_from_sa),
      .pb_dma_to_descriptor_memory_s1_waitrequest_from_sa                                     (pb_dma_to_descriptor_memory_s1_waitrequest_from_sa),
      .reset_n                                                                                (ddr3_top_phy_clk_out_reset_n),
      .sgdma_rx_descriptor_read_address                                                       (sgdma_rx_descriptor_read_address),
      .sgdma_rx_descriptor_read_address_to_slave                                              (sgdma_rx_descriptor_read_address_to_slave),
      .sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1                        (sgdma_rx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_latency_counter                                               (sgdma_rx_descriptor_read_latency_counter),
      .sgdma_rx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1              (sgdma_rx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_read                                                          (sgdma_rx_descriptor_read_read),
      .sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1                (sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register (sgdma_rx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register),
      .sgdma_rx_descriptor_read_readdata                                                      (sgdma_rx_descriptor_read_readdata),
      .sgdma_rx_descriptor_read_readdatavalid                                                 (sgdma_rx_descriptor_read_readdatavalid),
      .sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1                       (sgdma_rx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_waitrequest                                                   (sgdma_rx_descriptor_read_waitrequest)
    );

  sgdma_rx_descriptor_write_arbitrator the_sgdma_rx_descriptor_write
    (
      .clk                                                                        (ddr3_top_phy_clk_out),
      .d1_pb_dma_to_descriptor_memory_s1_end_xfer                                 (d1_pb_dma_to_descriptor_memory_s1_end_xfer),
      .pb_dma_to_descriptor_memory_s1_waitrequest_from_sa                         (pb_dma_to_descriptor_memory_s1_waitrequest_from_sa),
      .reset_n                                                                    (ddr3_top_phy_clk_out_reset_n),
      .sgdma_rx_descriptor_write_address                                          (sgdma_rx_descriptor_write_address),
      .sgdma_rx_descriptor_write_address_to_slave                                 (sgdma_rx_descriptor_write_address_to_slave),
      .sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1           (sgdma_rx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1 (sgdma_rx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1          (sgdma_rx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_waitrequest                                      (sgdma_rx_descriptor_write_waitrequest),
      .sgdma_rx_descriptor_write_write                                            (sgdma_rx_descriptor_write_write),
      .sgdma_rx_descriptor_write_writedata                                        (sgdma_rx_descriptor_write_writedata)
    );

  sgdma_rx_m_write_arbitrator the_sgdma_rx_m_write
    (
      .clk                                                      (ddr3_top_phy_clk_out),
      .d1_pb_dma_to_ddr3_top_s1_end_xfer                        (d1_pb_dma_to_ddr3_top_s1_end_xfer),
      .pb_dma_to_ddr3_top_s1_waitrequest_from_sa                (pb_dma_to_ddr3_top_s1_waitrequest_from_sa),
      .reset_n                                                  (ddr3_top_phy_clk_out_reset_n),
      .sgdma_rx_m_write_address                                 (sgdma_rx_m_write_address),
      .sgdma_rx_m_write_address_to_slave                        (sgdma_rx_m_write_address_to_slave),
      .sgdma_rx_m_write_byteenable                              (sgdma_rx_m_write_byteenable),
      .sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1           (sgdma_rx_m_write_granted_pb_dma_to_ddr3_top_s1),
      .sgdma_rx_m_write_qualified_request_pb_dma_to_ddr3_top_s1 (sgdma_rx_m_write_qualified_request_pb_dma_to_ddr3_top_s1),
      .sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1          (sgdma_rx_m_write_requests_pb_dma_to_ddr3_top_s1),
      .sgdma_rx_m_write_waitrequest                             (sgdma_rx_m_write_waitrequest),
      .sgdma_rx_m_write_write                                   (sgdma_rx_m_write_write),
      .sgdma_rx_m_write_writedata                               (sgdma_rx_m_write_writedata)
    );

  sgdma_rx the_sgdma_rx
    (
      .clk                           (ddr3_top_phy_clk_out),
      .csr_address                   (sgdma_rx_csr_address),
      .csr_chipselect                (sgdma_rx_csr_chipselect),
      .csr_irq                       (sgdma_rx_csr_irq),
      .csr_read                      (sgdma_rx_csr_read),
      .csr_readdata                  (sgdma_rx_csr_readdata),
      .csr_write                     (sgdma_rx_csr_write),
      .csr_writedata                 (sgdma_rx_csr_writedata),
      .descriptor_read_address       (sgdma_rx_descriptor_read_address),
      .descriptor_read_read          (sgdma_rx_descriptor_read_read),
      .descriptor_read_readdata      (sgdma_rx_descriptor_read_readdata),
      .descriptor_read_readdatavalid (sgdma_rx_descriptor_read_readdatavalid),
      .descriptor_read_waitrequest   (sgdma_rx_descriptor_read_waitrequest),
      .descriptor_write_address      (sgdma_rx_descriptor_write_address),
      .descriptor_write_waitrequest  (sgdma_rx_descriptor_write_waitrequest),
      .descriptor_write_write        (sgdma_rx_descriptor_write_write),
      .descriptor_write_writedata    (sgdma_rx_descriptor_write_writedata),
      .in_data                       (sgdma_rx_in_data),
      .in_empty                      (sgdma_rx_in_empty),
      .in_endofpacket                (sgdma_rx_in_endofpacket),
      .in_error                      (sgdma_rx_in_error),
      .in_ready                      (sgdma_rx_in_ready),
      .in_startofpacket              (sgdma_rx_in_startofpacket),
      .in_valid                      (sgdma_rx_in_valid),
      .m_write_address               (sgdma_rx_m_write_address),
      .m_write_byteenable            (sgdma_rx_m_write_byteenable),
      .m_write_waitrequest           (sgdma_rx_m_write_waitrequest),
      .m_write_write                 (sgdma_rx_m_write_write),
      .m_write_writedata             (sgdma_rx_m_write_writedata),
      .system_reset_n                (sgdma_rx_csr_reset_n)
    );

  sgdma_tx_csr_arbitrator the_sgdma_tx_csr
    (
      .clk                                            (ddr3_top_phy_clk_out),
      .d1_sgdma_tx_csr_end_xfer                       (d1_sgdma_tx_csr_end_xfer),
      .pb_cpu_to_io_m1_address_to_slave               (pb_cpu_to_io_m1_address_to_slave),
      .pb_cpu_to_io_m1_burstcount                     (pb_cpu_to_io_m1_burstcount),
      .pb_cpu_to_io_m1_chipselect                     (pb_cpu_to_io_m1_chipselect),
      .pb_cpu_to_io_m1_granted_sgdma_tx_csr           (pb_cpu_to_io_m1_granted_sgdma_tx_csr),
      .pb_cpu_to_io_m1_latency_counter                (pb_cpu_to_io_m1_latency_counter),
      .pb_cpu_to_io_m1_qualified_request_sgdma_tx_csr (pb_cpu_to_io_m1_qualified_request_sgdma_tx_csr),
      .pb_cpu_to_io_m1_read                           (pb_cpu_to_io_m1_read),
      .pb_cpu_to_io_m1_read_data_valid_sgdma_tx_csr   (pb_cpu_to_io_m1_read_data_valid_sgdma_tx_csr),
      .pb_cpu_to_io_m1_requests_sgdma_tx_csr          (pb_cpu_to_io_m1_requests_sgdma_tx_csr),
      .pb_cpu_to_io_m1_write                          (pb_cpu_to_io_m1_write),
      .pb_cpu_to_io_m1_writedata                      (pb_cpu_to_io_m1_writedata),
      .reset_n                                        (ddr3_top_phy_clk_out_reset_n),
      .sgdma_tx_csr_address                           (sgdma_tx_csr_address),
      .sgdma_tx_csr_chipselect                        (sgdma_tx_csr_chipselect),
      .sgdma_tx_csr_irq                               (sgdma_tx_csr_irq),
      .sgdma_tx_csr_irq_from_sa                       (sgdma_tx_csr_irq_from_sa),
      .sgdma_tx_csr_read                              (sgdma_tx_csr_read),
      .sgdma_tx_csr_readdata                          (sgdma_tx_csr_readdata),
      .sgdma_tx_csr_readdata_from_sa                  (sgdma_tx_csr_readdata_from_sa),
      .sgdma_tx_csr_reset_n                           (sgdma_tx_csr_reset_n),
      .sgdma_tx_csr_write                             (sgdma_tx_csr_write),
      .sgdma_tx_csr_writedata                         (sgdma_tx_csr_writedata)
    );

  sgdma_tx_descriptor_read_arbitrator the_sgdma_tx_descriptor_read
    (
      .clk                                                                                    (ddr3_top_phy_clk_out),
      .d1_pb_dma_to_descriptor_memory_s1_end_xfer                                             (d1_pb_dma_to_descriptor_memory_s1_end_xfer),
      .pb_dma_to_descriptor_memory_s1_readdata_from_sa                                        (pb_dma_to_descriptor_memory_s1_readdata_from_sa),
      .pb_dma_to_descriptor_memory_s1_waitrequest_from_sa                                     (pb_dma_to_descriptor_memory_s1_waitrequest_from_sa),
      .reset_n                                                                                (ddr3_top_phy_clk_out_reset_n),
      .sgdma_tx_descriptor_read_address                                                       (sgdma_tx_descriptor_read_address),
      .sgdma_tx_descriptor_read_address_to_slave                                              (sgdma_tx_descriptor_read_address_to_slave),
      .sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1                        (sgdma_tx_descriptor_read_granted_pb_dma_to_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_latency_counter                                               (sgdma_tx_descriptor_read_latency_counter),
      .sgdma_tx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1              (sgdma_tx_descriptor_read_qualified_request_pb_dma_to_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_read                                                          (sgdma_tx_descriptor_read_read),
      .sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1                (sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register (sgdma_tx_descriptor_read_read_data_valid_pb_dma_to_descriptor_memory_s1_shift_register),
      .sgdma_tx_descriptor_read_readdata                                                      (sgdma_tx_descriptor_read_readdata),
      .sgdma_tx_descriptor_read_readdatavalid                                                 (sgdma_tx_descriptor_read_readdatavalid),
      .sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1                       (sgdma_tx_descriptor_read_requests_pb_dma_to_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_waitrequest                                                   (sgdma_tx_descriptor_read_waitrequest)
    );

  sgdma_tx_descriptor_write_arbitrator the_sgdma_tx_descriptor_write
    (
      .clk                                                                        (ddr3_top_phy_clk_out),
      .d1_pb_dma_to_descriptor_memory_s1_end_xfer                                 (d1_pb_dma_to_descriptor_memory_s1_end_xfer),
      .pb_dma_to_descriptor_memory_s1_waitrequest_from_sa                         (pb_dma_to_descriptor_memory_s1_waitrequest_from_sa),
      .reset_n                                                                    (ddr3_top_phy_clk_out_reset_n),
      .sgdma_tx_descriptor_write_address                                          (sgdma_tx_descriptor_write_address),
      .sgdma_tx_descriptor_write_address_to_slave                                 (sgdma_tx_descriptor_write_address_to_slave),
      .sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1           (sgdma_tx_descriptor_write_granted_pb_dma_to_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1 (sgdma_tx_descriptor_write_qualified_request_pb_dma_to_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1          (sgdma_tx_descriptor_write_requests_pb_dma_to_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_waitrequest                                      (sgdma_tx_descriptor_write_waitrequest),
      .sgdma_tx_descriptor_write_write                                            (sgdma_tx_descriptor_write_write),
      .sgdma_tx_descriptor_write_writedata                                        (sgdma_tx_descriptor_write_writedata)
    );

  sgdma_tx_m_read_arbitrator the_sgdma_tx_m_read
    (
      .clk                                                                  (ddr3_top_phy_clk_out),
      .d1_pb_dma_to_ddr3_top_s1_end_xfer                                    (d1_pb_dma_to_ddr3_top_s1_end_xfer),
      .pb_dma_to_ddr3_top_s1_readdata_from_sa                               (pb_dma_to_ddr3_top_s1_readdata_from_sa),
      .pb_dma_to_ddr3_top_s1_waitrequest_from_sa                            (pb_dma_to_ddr3_top_s1_waitrequest_from_sa),
      .reset_n                                                              (ddr3_top_phy_clk_out_reset_n),
      .sgdma_tx_m_read_address                                              (sgdma_tx_m_read_address),
      .sgdma_tx_m_read_address_to_slave                                     (sgdma_tx_m_read_address_to_slave),
      .sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1                        (sgdma_tx_m_read_granted_pb_dma_to_ddr3_top_s1),
      .sgdma_tx_m_read_latency_counter                                      (sgdma_tx_m_read_latency_counter),
      .sgdma_tx_m_read_qualified_request_pb_dma_to_ddr3_top_s1              (sgdma_tx_m_read_qualified_request_pb_dma_to_ddr3_top_s1),
      .sgdma_tx_m_read_read                                                 (sgdma_tx_m_read_read),
      .sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1                (sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1),
      .sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1_shift_register (sgdma_tx_m_read_read_data_valid_pb_dma_to_ddr3_top_s1_shift_register),
      .sgdma_tx_m_read_readdata                                             (sgdma_tx_m_read_readdata),
      .sgdma_tx_m_read_readdatavalid                                        (sgdma_tx_m_read_readdatavalid),
      .sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1                       (sgdma_tx_m_read_requests_pb_dma_to_ddr3_top_s1),
      .sgdma_tx_m_read_waitrequest                                          (sgdma_tx_m_read_waitrequest)
    );

  sgdma_tx_out_arbitrator the_sgdma_tx_out
    (
      .clk                            (ddr3_top_phy_clk_out),
      .reset_n                        (ddr3_top_phy_clk_out_reset_n),
      .sgdma_tx_out_data              (sgdma_tx_out_data),
      .sgdma_tx_out_empty             (sgdma_tx_out_empty),
      .sgdma_tx_out_endofpacket       (sgdma_tx_out_endofpacket),
      .sgdma_tx_out_error             (sgdma_tx_out_error),
      .sgdma_tx_out_ready             (sgdma_tx_out_ready),
      .sgdma_tx_out_startofpacket     (sgdma_tx_out_startofpacket),
      .sgdma_tx_out_valid             (sgdma_tx_out_valid),
      .tse_mac_transmit_ready_from_sa (tse_mac_transmit_ready_from_sa)
    );

  sgdma_tx the_sgdma_tx
    (
      .clk                           (ddr3_top_phy_clk_out),
      .csr_address                   (sgdma_tx_csr_address),
      .csr_chipselect                (sgdma_tx_csr_chipselect),
      .csr_irq                       (sgdma_tx_csr_irq),
      .csr_read                      (sgdma_tx_csr_read),
      .csr_readdata                  (sgdma_tx_csr_readdata),
      .csr_write                     (sgdma_tx_csr_write),
      .csr_writedata                 (sgdma_tx_csr_writedata),
      .descriptor_read_address       (sgdma_tx_descriptor_read_address),
      .descriptor_read_read          (sgdma_tx_descriptor_read_read),
      .descriptor_read_readdata      (sgdma_tx_descriptor_read_readdata),
      .descriptor_read_readdatavalid (sgdma_tx_descriptor_read_readdatavalid),
      .descriptor_read_waitrequest   (sgdma_tx_descriptor_read_waitrequest),
      .descriptor_write_address      (sgdma_tx_descriptor_write_address),
      .descriptor_write_waitrequest  (sgdma_tx_descriptor_write_waitrequest),
      .descriptor_write_write        (sgdma_tx_descriptor_write_write),
      .descriptor_write_writedata    (sgdma_tx_descriptor_write_writedata),
      .m_read_address                (sgdma_tx_m_read_address),
      .m_read_read                   (sgdma_tx_m_read_read),
      .m_read_readdata               (sgdma_tx_m_read_readdata),
      .m_read_readdatavalid          (sgdma_tx_m_read_readdatavalid),
      .m_read_waitrequest            (sgdma_tx_m_read_waitrequest),
      .out_data                      (sgdma_tx_out_data),
      .out_empty                     (sgdma_tx_out_empty),
      .out_endofpacket               (sgdma_tx_out_endofpacket),
      .out_error                     (sgdma_tx_out_error),
      .out_ready                     (sgdma_tx_out_ready),
      .out_startofpacket             (sgdma_tx_out_startofpacket),
      .out_valid                     (sgdma_tx_out_valid),
      .system_reset_n                (sgdma_tx_csr_reset_n)
    );

  sysid_control_slave_arbitrator the_sysid_control_slave
    (
      .clk                                                   (ddr3_top_phy_clk_out),
      .d1_sysid_control_slave_end_xfer                       (d1_sysid_control_slave_end_xfer),
      .pb_cpu_to_io_m1_address_to_slave                      (pb_cpu_to_io_m1_address_to_slave),
      .pb_cpu_to_io_m1_burstcount                            (pb_cpu_to_io_m1_burstcount),
      .pb_cpu_to_io_m1_chipselect                            (pb_cpu_to_io_m1_chipselect),
      .pb_cpu_to_io_m1_granted_sysid_control_slave           (pb_cpu_to_io_m1_granted_sysid_control_slave),
      .pb_cpu_to_io_m1_latency_counter                       (pb_cpu_to_io_m1_latency_counter),
      .pb_cpu_to_io_m1_qualified_request_sysid_control_slave (pb_cpu_to_io_m1_qualified_request_sysid_control_slave),
      .pb_cpu_to_io_m1_read                                  (pb_cpu_to_io_m1_read),
      .pb_cpu_to_io_m1_read_data_valid_sysid_control_slave   (pb_cpu_to_io_m1_read_data_valid_sysid_control_slave),
      .pb_cpu_to_io_m1_requests_sysid_control_slave          (pb_cpu_to_io_m1_requests_sysid_control_slave),
      .pb_cpu_to_io_m1_write                                 (pb_cpu_to_io_m1_write),
      .reset_n                                               (ddr3_top_phy_clk_out_reset_n),
      .sysid_control_slave_address                           (sysid_control_slave_address),
      .sysid_control_slave_readdata                          (sysid_control_slave_readdata),
      .sysid_control_slave_readdata_from_sa                  (sysid_control_slave_readdata_from_sa),
      .sysid_control_slave_reset_n                           (sysid_control_slave_reset_n)
    );

  sysid the_sysid
    (
      .address  (sysid_control_slave_address),
      .clock    (sysid_control_slave_clock),
      .readdata (sysid_control_slave_readdata),
      .reset_n  (sysid_control_slave_reset_n)
    );

  tb_fsm_avalon_slave_arbitrator the_tb_fsm_avalon_slave
    (
      .clk                                               (ddr3_top_phy_clk_out),
      .d1_tb_fsm_avalon_slave_end_xfer                   (d1_tb_fsm_avalon_slave_end_xfer),
      .ext_flash_1_s1_wait_counter_eq_0                  (ext_flash_1_s1_wait_counter_eq_0),
      .ext_flash_s1_wait_counter_eq_0                    (ext_flash_s1_wait_counter_eq_0),
      .incoming_tb_fsm_data_with_Xs_converted_to_0       (incoming_tb_fsm_data_with_Xs_converted_to_0),
      .pb_cpu_to_fsm_m1_address_to_slave                 (pb_cpu_to_fsm_m1_address_to_slave),
      .pb_cpu_to_fsm_m1_burstcount                       (pb_cpu_to_fsm_m1_burstcount),
      .pb_cpu_to_fsm_m1_byteenable                       (pb_cpu_to_fsm_m1_byteenable),
      .pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1        (pb_cpu_to_fsm_m1_byteenable_ext_flash_1_s1),
      .pb_cpu_to_fsm_m1_byteenable_ext_flash_s1          (pb_cpu_to_fsm_m1_byteenable_ext_flash_s1),
      .pb_cpu_to_fsm_m1_chipselect                       (pb_cpu_to_fsm_m1_chipselect),
      .pb_cpu_to_fsm_m1_dbs_address                      (pb_cpu_to_fsm_m1_dbs_address),
      .pb_cpu_to_fsm_m1_dbs_write_16                     (pb_cpu_to_fsm_m1_dbs_write_16),
      .pb_cpu_to_fsm_m1_granted_ext_flash_1_s1           (pb_cpu_to_fsm_m1_granted_ext_flash_1_s1),
      .pb_cpu_to_fsm_m1_granted_ext_flash_s1             (pb_cpu_to_fsm_m1_granted_ext_flash_s1),
      .pb_cpu_to_fsm_m1_latency_counter                  (pb_cpu_to_fsm_m1_latency_counter),
      .pb_cpu_to_fsm_m1_qualified_request_ext_flash_1_s1 (pb_cpu_to_fsm_m1_qualified_request_ext_flash_1_s1),
      .pb_cpu_to_fsm_m1_qualified_request_ext_flash_s1   (pb_cpu_to_fsm_m1_qualified_request_ext_flash_s1),
      .pb_cpu_to_fsm_m1_read                             (pb_cpu_to_fsm_m1_read),
      .pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1   (pb_cpu_to_fsm_m1_read_data_valid_ext_flash_1_s1),
      .pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1     (pb_cpu_to_fsm_m1_read_data_valid_ext_flash_s1),
      .pb_cpu_to_fsm_m1_requests_ext_flash_1_s1          (pb_cpu_to_fsm_m1_requests_ext_flash_1_s1),
      .pb_cpu_to_fsm_m1_requests_ext_flash_s1            (pb_cpu_to_fsm_m1_requests_ext_flash_s1),
      .pb_cpu_to_fsm_m1_write                            (pb_cpu_to_fsm_m1_write),
      .reset_n                                           (ddr3_top_phy_clk_out_reset_n),
      .select_n_to_the_ext_flash                         (select_n_to_the_ext_flash),
      .select_n_to_the_ext_flash_1                       (select_n_to_the_ext_flash_1),
      .tb_fsm_address                                    (tb_fsm_address),
      .tb_fsm_data                                       (tb_fsm_data),
      .tb_fsm_readn                                      (tb_fsm_readn),
      .tb_fsm_writen                                     (tb_fsm_writen)
    );

  timer_1ms_s1_arbitrator the_timer_1ms_s1
    (
      .clk                                            (ddr3_top_phy_clk_out),
      .d1_timer_1ms_s1_end_xfer                       (d1_timer_1ms_s1_end_xfer),
      .pb_cpu_to_io_m1_address_to_slave               (pb_cpu_to_io_m1_address_to_slave),
      .pb_cpu_to_io_m1_burstcount                     (pb_cpu_to_io_m1_burstcount),
      .pb_cpu_to_io_m1_chipselect                     (pb_cpu_to_io_m1_chipselect),
      .pb_cpu_to_io_m1_granted_timer_1ms_s1           (pb_cpu_to_io_m1_granted_timer_1ms_s1),
      .pb_cpu_to_io_m1_latency_counter                (pb_cpu_to_io_m1_latency_counter),
      .pb_cpu_to_io_m1_qualified_request_timer_1ms_s1 (pb_cpu_to_io_m1_qualified_request_timer_1ms_s1),
      .pb_cpu_to_io_m1_read                           (pb_cpu_to_io_m1_read),
      .pb_cpu_to_io_m1_read_data_valid_timer_1ms_s1   (pb_cpu_to_io_m1_read_data_valid_timer_1ms_s1),
      .pb_cpu_to_io_m1_requests_timer_1ms_s1          (pb_cpu_to_io_m1_requests_timer_1ms_s1),
      .pb_cpu_to_io_m1_write                          (pb_cpu_to_io_m1_write),
      .pb_cpu_to_io_m1_writedata                      (pb_cpu_to_io_m1_writedata),
      .reset_n                                        (ddr3_top_phy_clk_out_reset_n),
      .timer_1ms_s1_address                           (timer_1ms_s1_address),
      .timer_1ms_s1_chipselect                        (timer_1ms_s1_chipselect),
      .timer_1ms_s1_irq                               (timer_1ms_s1_irq),
      .timer_1ms_s1_irq_from_sa                       (timer_1ms_s1_irq_from_sa),
      .timer_1ms_s1_readdata                          (timer_1ms_s1_readdata),
      .timer_1ms_s1_readdata_from_sa                  (timer_1ms_s1_readdata_from_sa),
      .timer_1ms_s1_reset_n                           (timer_1ms_s1_reset_n),
      .timer_1ms_s1_write_n                           (timer_1ms_s1_write_n),
      .timer_1ms_s1_writedata                         (timer_1ms_s1_writedata)
    );

  timer_1ms the_timer_1ms
    (
      .address    (timer_1ms_s1_address),
      .chipselect (timer_1ms_s1_chipselect),
      .clk        (ddr3_top_phy_clk_out),
      .irq        (timer_1ms_s1_irq),
      .readdata   (timer_1ms_s1_readdata),
      .reset_n    (timer_1ms_s1_reset_n),
      .write_n    (timer_1ms_s1_write_n),
      .writedata  (timer_1ms_s1_writedata)
    );

  tlb_miss_ram_1k_s1_arbitrator the_tlb_miss_ram_1k_s1
    (
      .clk                                                                           (ddr3_top_phy_clk_out),
      .cpu_tightly_coupled_instruction_master_0_address_to_slave                     (cpu_tightly_coupled_instruction_master_0_address_to_slave),
      .cpu_tightly_coupled_instruction_master_0_clken                                (cpu_tightly_coupled_instruction_master_0_clken),
      .cpu_tightly_coupled_instruction_master_0_granted_tlb_miss_ram_1k_s1           (cpu_tightly_coupled_instruction_master_0_granted_tlb_miss_ram_1k_s1),
      .cpu_tightly_coupled_instruction_master_0_latency_counter                      (cpu_tightly_coupled_instruction_master_0_latency_counter),
      .cpu_tightly_coupled_instruction_master_0_qualified_request_tlb_miss_ram_1k_s1 (cpu_tightly_coupled_instruction_master_0_qualified_request_tlb_miss_ram_1k_s1),
      .cpu_tightly_coupled_instruction_master_0_read                                 (cpu_tightly_coupled_instruction_master_0_read),
      .cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1   (cpu_tightly_coupled_instruction_master_0_read_data_valid_tlb_miss_ram_1k_s1),
      .cpu_tightly_coupled_instruction_master_0_requests_tlb_miss_ram_1k_s1          (cpu_tightly_coupled_instruction_master_0_requests_tlb_miss_ram_1k_s1),
      .d1_tlb_miss_ram_1k_s1_end_xfer                                                (d1_tlb_miss_ram_1k_s1_end_xfer),
      .reset_n                                                                       (ddr3_top_phy_clk_out_reset_n),
      .tlb_miss_ram_1k_s1_address                                                    (tlb_miss_ram_1k_s1_address),
      .tlb_miss_ram_1k_s1_byteenable                                                 (tlb_miss_ram_1k_s1_byteenable),
      .tlb_miss_ram_1k_s1_chipselect                                                 (tlb_miss_ram_1k_s1_chipselect),
      .tlb_miss_ram_1k_s1_clken                                                      (tlb_miss_ram_1k_s1_clken),
      .tlb_miss_ram_1k_s1_readdata                                                   (tlb_miss_ram_1k_s1_readdata),
      .tlb_miss_ram_1k_s1_readdata_from_sa                                           (tlb_miss_ram_1k_s1_readdata_from_sa),
      .tlb_miss_ram_1k_s1_reset                                                      (tlb_miss_ram_1k_s1_reset),
      .tlb_miss_ram_1k_s1_write                                                      (tlb_miss_ram_1k_s1_write),
      .tlb_miss_ram_1k_s1_writedata                                                  (tlb_miss_ram_1k_s1_writedata)
    );

  tlb_miss_ram_1k_s2_arbitrator the_tlb_miss_ram_1k_s2
    (
      .clk                                                                    (ddr3_top_phy_clk_out),
      .cpu_tightly_coupled_data_master_0_address_to_slave                     (cpu_tightly_coupled_data_master_0_address_to_slave),
      .cpu_tightly_coupled_data_master_0_byteenable                           (cpu_tightly_coupled_data_master_0_byteenable),
      .cpu_tightly_coupled_data_master_0_clken                                (cpu_tightly_coupled_data_master_0_clken),
      .cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2           (cpu_tightly_coupled_data_master_0_granted_tlb_miss_ram_1k_s2),
      .cpu_tightly_coupled_data_master_0_latency_counter                      (cpu_tightly_coupled_data_master_0_latency_counter),
      .cpu_tightly_coupled_data_master_0_qualified_request_tlb_miss_ram_1k_s2 (cpu_tightly_coupled_data_master_0_qualified_request_tlb_miss_ram_1k_s2),
      .cpu_tightly_coupled_data_master_0_read                                 (cpu_tightly_coupled_data_master_0_read),
      .cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2   (cpu_tightly_coupled_data_master_0_read_data_valid_tlb_miss_ram_1k_s2),
      .cpu_tightly_coupled_data_master_0_requests_tlb_miss_ram_1k_s2          (cpu_tightly_coupled_data_master_0_requests_tlb_miss_ram_1k_s2),
      .cpu_tightly_coupled_data_master_0_write                                (cpu_tightly_coupled_data_master_0_write),
      .cpu_tightly_coupled_data_master_0_writedata                            (cpu_tightly_coupled_data_master_0_writedata),
      .d1_tlb_miss_ram_1k_s2_end_xfer                                         (d1_tlb_miss_ram_1k_s2_end_xfer),
      .reset_n                                                                (ddr3_top_phy_clk_out_reset_n),
      .tlb_miss_ram_1k_s2_address                                             (tlb_miss_ram_1k_s2_address),
      .tlb_miss_ram_1k_s2_byteenable                                          (tlb_miss_ram_1k_s2_byteenable),
      .tlb_miss_ram_1k_s2_chipselect                                          (tlb_miss_ram_1k_s2_chipselect),
      .tlb_miss_ram_1k_s2_clken                                               (tlb_miss_ram_1k_s2_clken),
      .tlb_miss_ram_1k_s2_readdata                                            (tlb_miss_ram_1k_s2_readdata),
      .tlb_miss_ram_1k_s2_readdata_from_sa                                    (tlb_miss_ram_1k_s2_readdata_from_sa),
      .tlb_miss_ram_1k_s2_reset                                               (tlb_miss_ram_1k_s2_reset),
      .tlb_miss_ram_1k_s2_write                                               (tlb_miss_ram_1k_s2_write),
      .tlb_miss_ram_1k_s2_writedata                                           (tlb_miss_ram_1k_s2_writedata)
    );

  tlb_miss_ram_1k the_tlb_miss_ram_1k
    (
      .address     (tlb_miss_ram_1k_s1_address),
      .address2    (tlb_miss_ram_1k_s2_address),
      .byteenable  (tlb_miss_ram_1k_s1_byteenable),
      .byteenable2 (tlb_miss_ram_1k_s2_byteenable),
      .chipselect  (tlb_miss_ram_1k_s1_chipselect),
      .chipselect2 (tlb_miss_ram_1k_s2_chipselect),
      .clk         (ddr3_top_phy_clk_out),
      .clk2        (ddr3_top_phy_clk_out),
      .clken       (tlb_miss_ram_1k_s1_clken),
      .clken2      (tlb_miss_ram_1k_s2_clken),
      .readdata    (tlb_miss_ram_1k_s1_readdata),
      .readdata2   (tlb_miss_ram_1k_s2_readdata),
      .reset       (tlb_miss_ram_1k_s1_reset),
      .reset2      (tlb_miss_ram_1k_s2_reset),
      .write       (tlb_miss_ram_1k_s1_write),
      .write2      (tlb_miss_ram_1k_s2_write),
      .writedata   (tlb_miss_ram_1k_s1_writedata),
      .writedata2  (tlb_miss_ram_1k_s2_writedata)
    );

  tse_mac_control_port_arbitrator the_tse_mac_control_port
    (
      .clk                                                    (ddr3_top_phy_clk_out),
      .d1_tse_mac_control_port_end_xfer                       (d1_tse_mac_control_port_end_xfer),
      .pb_cpu_to_io_m1_address_to_slave                       (pb_cpu_to_io_m1_address_to_slave),
      .pb_cpu_to_io_m1_burstcount                             (pb_cpu_to_io_m1_burstcount),
      .pb_cpu_to_io_m1_chipselect                             (pb_cpu_to_io_m1_chipselect),
      .pb_cpu_to_io_m1_granted_tse_mac_control_port           (pb_cpu_to_io_m1_granted_tse_mac_control_port),
      .pb_cpu_to_io_m1_latency_counter                        (pb_cpu_to_io_m1_latency_counter),
      .pb_cpu_to_io_m1_qualified_request_tse_mac_control_port (pb_cpu_to_io_m1_qualified_request_tse_mac_control_port),
      .pb_cpu_to_io_m1_read                                   (pb_cpu_to_io_m1_read),
      .pb_cpu_to_io_m1_read_data_valid_tse_mac_control_port   (pb_cpu_to_io_m1_read_data_valid_tse_mac_control_port),
      .pb_cpu_to_io_m1_requests_tse_mac_control_port          (pb_cpu_to_io_m1_requests_tse_mac_control_port),
      .pb_cpu_to_io_m1_write                                  (pb_cpu_to_io_m1_write),
      .pb_cpu_to_io_m1_writedata                              (pb_cpu_to_io_m1_writedata),
      .reset_n                                                (ddr3_top_phy_clk_out_reset_n),
      .tse_mac_control_port_address                           (tse_mac_control_port_address),
      .tse_mac_control_port_read                              (tse_mac_control_port_read),
      .tse_mac_control_port_readdata                          (tse_mac_control_port_readdata),
      .tse_mac_control_port_readdata_from_sa                  (tse_mac_control_port_readdata_from_sa),
      .tse_mac_control_port_reset                             (tse_mac_control_port_reset),
      .tse_mac_control_port_waitrequest                       (tse_mac_control_port_waitrequest),
      .tse_mac_control_port_waitrequest_from_sa               (tse_mac_control_port_waitrequest_from_sa),
      .tse_mac_control_port_write                             (tse_mac_control_port_write),
      .tse_mac_control_port_writedata                         (tse_mac_control_port_writedata)
    );

  tse_mac_transmit_arbitrator the_tse_mac_transmit
    (
      .clk                            (ddr3_top_phy_clk_out),
      .reset_n                        (ddr3_top_phy_clk_out_reset_n),
      .sgdma_tx_out_data              (sgdma_tx_out_data),
      .sgdma_tx_out_empty             (sgdma_tx_out_empty),
      .sgdma_tx_out_endofpacket       (sgdma_tx_out_endofpacket),
      .sgdma_tx_out_error             (sgdma_tx_out_error),
      .sgdma_tx_out_startofpacket     (sgdma_tx_out_startofpacket),
      .sgdma_tx_out_valid             (sgdma_tx_out_valid),
      .tse_mac_transmit_data          (tse_mac_transmit_data),
      .tse_mac_transmit_empty         (tse_mac_transmit_empty),
      .tse_mac_transmit_endofpacket   (tse_mac_transmit_endofpacket),
      .tse_mac_transmit_error         (tse_mac_transmit_error),
      .tse_mac_transmit_ready         (tse_mac_transmit_ready),
      .tse_mac_transmit_ready_from_sa (tse_mac_transmit_ready_from_sa),
      .tse_mac_transmit_startofpacket (tse_mac_transmit_startofpacket),
      .tse_mac_transmit_valid         (tse_mac_transmit_valid)
    );

  tse_mac_receive_arbitrator the_tse_mac_receive
    (
      .clk                           (ddr3_top_phy_clk_out),
      .reset_n                       (ddr3_top_phy_clk_out_reset_n),
      .sgdma_rx_in_ready_from_sa     (sgdma_rx_in_ready_from_sa),
      .tse_mac_receive_data          (tse_mac_receive_data),
      .tse_mac_receive_empty         (tse_mac_receive_empty),
      .tse_mac_receive_endofpacket   (tse_mac_receive_endofpacket),
      .tse_mac_receive_error         (tse_mac_receive_error),
      .tse_mac_receive_ready         (tse_mac_receive_ready),
      .tse_mac_receive_startofpacket (tse_mac_receive_startofpacket),
      .tse_mac_receive_valid         (tse_mac_receive_valid)
    );

  tse_mac the_tse_mac
    (
      .address        (tse_mac_control_port_address),
      .clk            (ddr3_top_phy_clk_out),
      .ff_rx_clk      (ddr3_top_phy_clk_out),
      .ff_rx_data     (tse_mac_receive_data),
      .ff_rx_dval     (tse_mac_receive_valid),
      .ff_rx_eop      (tse_mac_receive_endofpacket),
      .ff_rx_mod      (tse_mac_receive_empty),
      .ff_rx_rdy      (tse_mac_receive_ready),
      .ff_rx_sop      (tse_mac_receive_startofpacket),
      .ff_tx_clk      (ddr3_top_phy_clk_out),
      .ff_tx_data     (tse_mac_transmit_data),
      .ff_tx_eop      (tse_mac_transmit_endofpacket),
      .ff_tx_err      (tse_mac_transmit_error),
      .ff_tx_mod      (tse_mac_transmit_empty),
      .ff_tx_rdy      (tse_mac_transmit_ready),
      .ff_tx_sop      (tse_mac_transmit_startofpacket),
      .ff_tx_wren     (tse_mac_transmit_valid),
      .led_an         (led_an_from_the_tse_mac),
      .led_char_err   (led_char_err_from_the_tse_mac),
      .led_col        (led_col_from_the_tse_mac),
      .led_crs        (led_crs_from_the_tse_mac),
      .led_disp_err   (led_disp_err_from_the_tse_mac),
      .led_link       (led_link_from_the_tse_mac),
      .mdc            (mdc_from_the_tse_mac),
      .mdio_in        (mdio_in_to_the_tse_mac),
      .mdio_oen       (mdio_oen_from_the_tse_mac),
      .mdio_out       (mdio_out_from_the_tse_mac),
      .read           (tse_mac_control_port_read),
      .readdata       (tse_mac_control_port_readdata),
      .ref_clk        (ref_clk_to_the_tse_mac),
      .reset          (tse_mac_control_port_reset),
      .rx_err         (tse_mac_receive_error),
      .rx_recovclkout (rx_recovclkout_from_the_tse_mac),
      .rxp            (rxp_to_the_tse_mac),
      .txp            (txp_from_the_tse_mac),
      .waitrequest    (tse_mac_control_port_waitrequest),
      .write          (tse_mac_control_port_write),
      .writedata      (tse_mac_control_port_writedata)
    );

  uart_s1_arbitrator the_uart_s1
    (
      .clk                                       (ddr3_top_phy_clk_out),
      .d1_uart_s1_end_xfer                       (d1_uart_s1_end_xfer),
      .pb_cpu_to_io_m1_address_to_slave          (pb_cpu_to_io_m1_address_to_slave),
      .pb_cpu_to_io_m1_burstcount                (pb_cpu_to_io_m1_burstcount),
      .pb_cpu_to_io_m1_chipselect                (pb_cpu_to_io_m1_chipselect),
      .pb_cpu_to_io_m1_granted_uart_s1           (pb_cpu_to_io_m1_granted_uart_s1),
      .pb_cpu_to_io_m1_latency_counter           (pb_cpu_to_io_m1_latency_counter),
      .pb_cpu_to_io_m1_qualified_request_uart_s1 (pb_cpu_to_io_m1_qualified_request_uart_s1),
      .pb_cpu_to_io_m1_read                      (pb_cpu_to_io_m1_read),
      .pb_cpu_to_io_m1_read_data_valid_uart_s1   (pb_cpu_to_io_m1_read_data_valid_uart_s1),
      .pb_cpu_to_io_m1_requests_uart_s1          (pb_cpu_to_io_m1_requests_uart_s1),
      .pb_cpu_to_io_m1_write                     (pb_cpu_to_io_m1_write),
      .pb_cpu_to_io_m1_writedata                 (pb_cpu_to_io_m1_writedata),
      .reset_n                                   (ddr3_top_phy_clk_out_reset_n),
      .uart_s1_address                           (uart_s1_address),
      .uart_s1_begintransfer                     (uart_s1_begintransfer),
      .uart_s1_chipselect                        (uart_s1_chipselect),
      .uart_s1_dataavailable                     (uart_s1_dataavailable),
      .uart_s1_dataavailable_from_sa             (uart_s1_dataavailable_from_sa),
      .uart_s1_irq                               (uart_s1_irq),
      .uart_s1_irq_from_sa                       (uart_s1_irq_from_sa),
      .uart_s1_read_n                            (uart_s1_read_n),
      .uart_s1_readdata                          (uart_s1_readdata),
      .uart_s1_readdata_from_sa                  (uart_s1_readdata_from_sa),
      .uart_s1_readyfordata                      (uart_s1_readyfordata),
      .uart_s1_readyfordata_from_sa              (uart_s1_readyfordata_from_sa),
      .uart_s1_reset_n                           (uart_s1_reset_n),
      .uart_s1_write_n                           (uart_s1_write_n),
      .uart_s1_writedata                         (uart_s1_writedata)
    );

  uart the_uart
    (
      .address       (uart_s1_address),
      .begintransfer (uart_s1_begintransfer),
      .chipselect    (uart_s1_chipselect),
      .clk           (ddr3_top_phy_clk_out),
      .dataavailable (uart_s1_dataavailable),
      .irq           (uart_s1_irq),
      .read_n        (uart_s1_read_n),
      .readdata      (uart_s1_readdata),
      .readyfordata  (uart_s1_readyfordata),
      .reset_n       (uart_s1_reset_n),
      .rxd           (rxd_to_the_uart),
      .txd           (txd_from_the_uart),
      .write_n       (uart_s1_write_n),
      .writedata     (uart_s1_writedata)
    );

  //reset is asserted asynchronously and deasserted synchronously
  ghrd_4sgx230_sopc_reset_ddr3_top_phy_clk_out_domain_synch_module ghrd_4sgx230_sopc_reset_ddr3_top_phy_clk_out_domain_synch
    (
      .clk      (ddr3_top_phy_clk_out),
      .data_in  (1'b1),
      .data_out (ddr3_top_phy_clk_out_reset_n),
      .reset_n  (reset_n_sources)
    );

  //pb_cpu_to_ddr3_top_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign pb_cpu_to_ddr3_top_m1_endofpacket = 0;

  //pb_cpu_to_fsm_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign pb_cpu_to_fsm_m1_endofpacket = 0;

  //pb_cpu_to_io_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign pb_cpu_to_io_m1_endofpacket = 0;

  //pb_dma_to_ddr3_top_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign pb_dma_to_ddr3_top_m1_endofpacket = 0;

  //pb_dma_to_descriptor_memory_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign pb_dma_to_descriptor_memory_m1_endofpacket = 0;

  //sysid_control_slave_clock of type clock does not connect to anything so wire it to default (0)
  assign sysid_control_slave_clock = 0;


endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_flash_lane0_module (
                                // inputs:
                                 data,
                                 rdaddress,
                                 rdclken,
                                 wraddress,
                                 wrclock,
                                 wren,

                                // outputs:
                                 q
                              )
;

  output  [  7: 0] q;
  input   [  7: 0] data;
  input   [ 23: 0] rdaddress;
  input            rdclken;
  input   [ 23: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [  7: 0] mem_array [16777215: 0];
  wire    [  7: 0] q;
  reg     [ 23: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      read_address = rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("ext_flash_lane0.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ext_flash_lane0.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 24,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_flash_lane1_module (
                                // inputs:
                                 data,
                                 rdaddress,
                                 rdclken,
                                 wraddress,
                                 wrclock,
                                 wren,

                                // outputs:
                                 q
                              )
;

  output  [  7: 0] q;
  input   [  7: 0] data;
  input   [ 23: 0] rdaddress;
  input            rdclken;
  input   [ 23: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [  7: 0] mem_array [16777215: 0];
  wire    [  7: 0] q;
  reg     [ 23: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      read_address = rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("ext_flash_lane1.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ext_flash_lane1.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 24,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_flash (
                   // inputs:
                    address,
                    read_n,
                    select_n,
                    write_n,

                   // outputs:
                    data
                 )
;

  inout   [ 15: 0] data;
  input   [ 23: 0] address;
  input            read_n;
  input            select_n;
  input            write_n;

  wire    [ 15: 0] data;
  wire    [  7: 0] data_0;
  wire    [  7: 0] data_1;
  wire    [ 15: 0] logic_vector_gasket;
  wire    [  7: 0] q_0;
  wire    [  7: 0] q_1;
  //s1, which is an e_ptf_slave

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  assign logic_vector_gasket = data;
  assign data_0 = logic_vector_gasket[7 : 0];
  //ext_flash_lane0, which is an e_ram
  ext_flash_lane0_module ext_flash_lane0
    (
      .data      (data_0),
      .q         (q_0),
      .rdaddress (address),
      .rdclken   (1'b1),
      .wraddress (address),
      .wrclock   (write_n),
      .wren      (~select_n)
    );

  assign data_1 = logic_vector_gasket[15 : 8];
  //ext_flash_lane1, which is an e_ram
  ext_flash_lane1_module ext_flash_lane1
    (
      .data      (data_1),
      .q         (q_1),
      .rdaddress (address),
      .rdclken   (1'b1),
      .wraddress (address),
      .wrclock   (write_n),
      .wren      (~select_n)
    );

  assign data = (~select_n & ~read_n)? {q_1,
    q_0}: {16{1'bz}};


//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_flash_1_lane0_module (
                                  // inputs:
                                   data,
                                   rdaddress,
                                   rdclken,
                                   wraddress,
                                   wrclock,
                                   wren,

                                  // outputs:
                                   q
                                )
;

  output  [  7: 0] q;
  input   [  7: 0] data;
  input   [ 23: 0] rdaddress;
  input            rdclken;
  input   [ 23: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [  7: 0] mem_array [16777215: 0];
  wire    [  7: 0] q;
  reg     [ 23: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      read_address = rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("ext_flash_1_lane0.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ext_flash_1_lane0.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 24,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_flash_1_lane1_module (
                                  // inputs:
                                   data,
                                   rdaddress,
                                   rdclken,
                                   wraddress,
                                   wrclock,
                                   wren,

                                  // outputs:
                                   q
                                )
;

  output  [  7: 0] q;
  input   [  7: 0] data;
  input   [ 23: 0] rdaddress;
  input            rdclken;
  input   [ 23: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [  7: 0] mem_array [16777215: 0];
  wire    [  7: 0] q;
  reg     [ 23: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      read_address = rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("ext_flash_1_lane1.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ext_flash_1_lane1.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 24,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_flash_1 (
                     // inputs:
                      address,
                      read_n,
                      select_n,
                      write_n,

                     // outputs:
                      data
                   )
;

  inout   [ 15: 0] data;
  input   [ 23: 0] address;
  input            read_n;
  input            select_n;
  input            write_n;

  wire    [ 15: 0] data;
  wire    [  7: 0] data_0;
  wire    [  7: 0] data_1;
  wire    [ 15: 0] logic_vector_gasket;
  wire    [  7: 0] q_0;
  wire    [  7: 0] q_1;
  //s1, which is an e_ptf_slave

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  assign logic_vector_gasket = data;
  assign data_0 = logic_vector_gasket[7 : 0];
  //ext_flash_1_lane0, which is an e_ram
  ext_flash_1_lane0_module ext_flash_1_lane0
    (
      .data      (data_0),
      .q         (q_0),
      .rdaddress (address),
      .rdclken   (1'b1),
      .wraddress (address),
      .wrclock   (write_n),
      .wren      (~select_n)
    );

  assign data_1 = logic_vector_gasket[15 : 8];
  //ext_flash_1_lane1, which is an e_ram
  ext_flash_1_lane1_module ext_flash_1_lane1
    (
      .data      (data_1),
      .q         (q_1),
      .rdaddress (address),
      .rdclken   (1'b1),
      .wraddress (address),
      .wrclock   (write_n),
      .wren      (~select_n)
    );

  assign data = (~select_n & ~read_n)? {q_1,
    q_0}: {16{1'bz}};


//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


//synthesis translate_off



// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE

// AND HERE WILL BE PRESERVED </ALTERA_NOTE>


// If user logic components use Altsync_Ram with convert_hex2ver.dll,
// set USE_convert_hex2ver in the user comments section above

// `ifdef USE_convert_hex2ver
// `else
// `define NO_PLI 1
// `endif

`include "/acds_builds/SJ/nightly/10.1/149/l32/acds/quartus/eda/sim_lib/altera_mf.v"
`include "/acds_builds/SJ/nightly/10.1/149/l32/acds/quartus/eda/sim_lib/220model.v"
`include "/acds_builds/SJ/nightly/10.1/149/l32/acds/quartus/eda/sim_lib/sgate.v"
`include "/acds_builds/SJ/nightly/10.1/149/l32/acds/quartus/eda/sim_lib/stratixiigx_hssi_atoms.v"
`include "/acds_builds/SJ/nightly/10.1/149/l32/acds/quartus/eda/sim_lib/stratixiv_hssi_atoms.v"
`include "tse_mac.vo"
`include "tse_mac_loopback.v"
`include "descriptor_memory.v"
`include "uart.v"
`include "sysid.v"
`include "button_pio.v"
`include "pb_cpu_to_io.v"
`include "led_pio.v"
`include "jtag_uart.v"
`include "tlb_miss_ram_1k.v"
`include "sgdma_rx.v"
`include "cpu_test_bench.v"
`include "cpu_mult_cell.v"
`include "cpu_oci_test_bench.v"
`include "cpu_jtag_debug_module_tck.v"
`include "cpu_jtag_debug_module_sysclk.v"
`include "cpu_jtag_debug_module_wrapper.v"
`include "cpu.v"
`include "pb_dma_to_ddr3_top.v"
`include "pb_cpu_to_fsm.v"
`include "pb_dma_to_descriptor_memory.v"
`include "sgdma_tx.v"
`include "pb_cpu_to_ddr3_top.v"
`include "timer_1ms.v"
`include "dipsw_pio.v"

`timescale 1ns / 1ps

module test_bench 
;


  wire             aux_scan_clk_from_the_ddr3_top;
  wire             aux_scan_clk_reset_n_from_the_ddr3_top;
  wire             clk;
  reg              clkin_100;
  wire             ddr3_top_aux_full_rate_clk_out;
  wire             ddr3_top_aux_half_rate_clk_out;
  wire             ddr3_top_phy_clk_out;
  wire             dll_reference_clk_from_the_ddr3_top;
  wire    [  5: 0] dqs_delay_ctrl_export_from_the_ddr3_top;
  wire             global_reset_n_to_the_ddr3_top;
  wire    [  2: 0] in_port_to_the_button_pio;
  wire    [  7: 0] in_port_to_the_dipsw_pio;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  wire             led_an_from_the_tse_mac;
  wire             led_char_err_from_the_tse_mac;
  wire             led_col_from_the_tse_mac;
  wire             led_crs_from_the_tse_mac;
  wire             led_disp_err_from_the_tse_mac;
  wire             led_link_from_the_tse_mac;
  wire             local_init_done_from_the_ddr3_top;
  wire             local_refresh_ack_from_the_ddr3_top;
  wire             local_wdata_req_from_the_ddr3_top;
  wire             mdc_from_the_tse_mac;
  wire             mdio_in_to_the_tse_mac;
  wire             mdio_oen_from_the_tse_mac;
  wire             mdio_out_from_the_tse_mac;
  wire    [ 12: 0] mem_addr_from_the_ddr3_top;
  wire    [  2: 0] mem_ba_from_the_ddr3_top;
  wire             mem_cas_n_from_the_ddr3_top;
  wire             mem_cke_from_the_ddr3_top;
  wire             mem_clk_n_to_and_from_the_ddr3_top;
  wire             mem_clk_to_and_from_the_ddr3_top;
  wire             mem_cs_n_from_the_ddr3_top;
  wire    [  1: 0] mem_dm_from_the_ddr3_top;
  wire    [ 15: 0] mem_dq_to_and_from_the_ddr3_top;
  wire    [  1: 0] mem_dqs_to_and_from_the_ddr3_top;
  wire    [  1: 0] mem_dqsn_to_and_from_the_ddr3_top;
  wire             mem_odt_from_the_ddr3_top;
  wire             mem_ras_n_from_the_ddr3_top;
  wire             mem_reset_n_from_the_ddr3_top;
  wire             mem_we_n_from_the_ddr3_top;
  wire    [ 13: 0] oct_ctl_rs_value_to_the_ddr3_top;
  wire    [ 13: 0] oct_ctl_rt_value_to_the_ddr3_top;
  wire    [ 15: 0] out_port_from_the_led_pio;
  wire             pb_cpu_to_ddr3_top_m1_debugaccess;
  wire             pb_cpu_to_ddr3_top_m1_endofpacket;
  wire             pb_cpu_to_ddr3_top_s1_endofpacket_from_sa;
  wire             pb_cpu_to_fsm_m1_debugaccess;
  wire             pb_cpu_to_fsm_m1_endofpacket;
  wire             pb_cpu_to_fsm_s1_endofpacket_from_sa;
  wire             pb_cpu_to_io_m1_debugaccess;
  wire             pb_cpu_to_io_m1_endofpacket;
  wire             pb_cpu_to_io_s1_endofpacket_from_sa;
  wire             pb_dma_to_ddr3_top_m1_debugaccess;
  wire             pb_dma_to_ddr3_top_m1_endofpacket;
  wire             pb_dma_to_ddr3_top_s1_endofpacket_from_sa;
  wire             pb_dma_to_descriptor_memory_m1_debugaccess;
  wire             pb_dma_to_descriptor_memory_m1_endofpacket;
  wire             pb_dma_to_descriptor_memory_s1_endofpacket_from_sa;
  wire             ref_clk_to_the_tse_mac;
  reg              reset_n;
  wire             reset_phy_clk_n_from_the_ddr3_top;
  wire             rx_recovclkout_from_the_tse_mac;
  wire             rxd_to_the_uart;
  wire             rxp_to_the_tse_mac;
  wire             select_n_to_the_ext_flash;
  wire             select_n_to_the_ext_flash_1;
  wire             sysid_control_slave_clock;
  wire    [ 24: 0] tb_fsm_address;
  wire    [ 15: 0] tb_fsm_data;
  wire             tb_fsm_readn;
  wire             tb_fsm_writen;
  wire             txd_from_the_uart;
  wire             txp_from_the_tse_mac;
  wire             uart_s1_dataavailable_from_sa;
  wire             uart_s1_readyfordata_from_sa;


// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
//  add your signals and additional architecture here
// AND HERE WILL BE PRESERVED </ALTERA_NOTE>

  //Set us up the Dut
  ghrd_4sgx230_sopc DUT
    (
      .aux_scan_clk_from_the_ddr3_top          (aux_scan_clk_from_the_ddr3_top),
      .aux_scan_clk_reset_n_from_the_ddr3_top  (aux_scan_clk_reset_n_from_the_ddr3_top),
      .clkin_100                               (clkin_100),
      .ddr3_top_aux_full_rate_clk_out          (ddr3_top_aux_full_rate_clk_out),
      .ddr3_top_aux_half_rate_clk_out          (ddr3_top_aux_half_rate_clk_out),
      .ddr3_top_phy_clk_out                    (ddr3_top_phy_clk_out),
      .dll_reference_clk_from_the_ddr3_top     (dll_reference_clk_from_the_ddr3_top),
      .dqs_delay_ctrl_export_from_the_ddr3_top (dqs_delay_ctrl_export_from_the_ddr3_top),
      .global_reset_n_to_the_ddr3_top          (global_reset_n_to_the_ddr3_top),
      .in_port_to_the_button_pio               (in_port_to_the_button_pio),
      .in_port_to_the_dipsw_pio                (in_port_to_the_dipsw_pio),
      .led_an_from_the_tse_mac                 (led_an_from_the_tse_mac),
      .led_char_err_from_the_tse_mac           (led_char_err_from_the_tse_mac),
      .led_col_from_the_tse_mac                (led_col_from_the_tse_mac),
      .led_crs_from_the_tse_mac                (led_crs_from_the_tse_mac),
      .led_disp_err_from_the_tse_mac           (led_disp_err_from_the_tse_mac),
      .led_link_from_the_tse_mac               (led_link_from_the_tse_mac),
      .local_init_done_from_the_ddr3_top       (local_init_done_from_the_ddr3_top),
      .local_refresh_ack_from_the_ddr3_top     (local_refresh_ack_from_the_ddr3_top),
      .local_wdata_req_from_the_ddr3_top       (local_wdata_req_from_the_ddr3_top),
      .mdc_from_the_tse_mac                    (mdc_from_the_tse_mac),
      .mdio_in_to_the_tse_mac                  (mdio_in_to_the_tse_mac),
      .mdio_oen_from_the_tse_mac               (mdio_oen_from_the_tse_mac),
      .mdio_out_from_the_tse_mac               (mdio_out_from_the_tse_mac),
      .mem_addr_from_the_ddr3_top              (mem_addr_from_the_ddr3_top),
      .mem_ba_from_the_ddr3_top                (mem_ba_from_the_ddr3_top),
      .mem_cas_n_from_the_ddr3_top             (mem_cas_n_from_the_ddr3_top),
      .mem_cke_from_the_ddr3_top               (mem_cke_from_the_ddr3_top),
      .mem_clk_n_to_and_from_the_ddr3_top      (mem_clk_n_to_and_from_the_ddr3_top),
      .mem_clk_to_and_from_the_ddr3_top        (mem_clk_to_and_from_the_ddr3_top),
      .mem_cs_n_from_the_ddr3_top              (mem_cs_n_from_the_ddr3_top),
      .mem_dm_from_the_ddr3_top                (mem_dm_from_the_ddr3_top),
      .mem_dq_to_and_from_the_ddr3_top         (mem_dq_to_and_from_the_ddr3_top),
      .mem_dqs_to_and_from_the_ddr3_top        (mem_dqs_to_and_from_the_ddr3_top),
      .mem_dqsn_to_and_from_the_ddr3_top       (mem_dqsn_to_and_from_the_ddr3_top),
      .mem_odt_from_the_ddr3_top               (mem_odt_from_the_ddr3_top),
      .mem_ras_n_from_the_ddr3_top             (mem_ras_n_from_the_ddr3_top),
      .mem_reset_n_from_the_ddr3_top           (mem_reset_n_from_the_ddr3_top),
      .mem_we_n_from_the_ddr3_top              (mem_we_n_from_the_ddr3_top),
      .oct_ctl_rs_value_to_the_ddr3_top        (oct_ctl_rs_value_to_the_ddr3_top),
      .oct_ctl_rt_value_to_the_ddr3_top        (oct_ctl_rt_value_to_the_ddr3_top),
      .out_port_from_the_led_pio               (out_port_from_the_led_pio),
      .ref_clk_to_the_tse_mac                  (ref_clk_to_the_tse_mac),
      .reset_n                                 (reset_n),
      .reset_phy_clk_n_from_the_ddr3_top       (reset_phy_clk_n_from_the_ddr3_top),
      .rx_recovclkout_from_the_tse_mac         (rx_recovclkout_from_the_tse_mac),
      .rxd_to_the_uart                         (rxd_to_the_uart),
      .rxp_to_the_tse_mac                      (rxp_to_the_tse_mac),
      .select_n_to_the_ext_flash               (select_n_to_the_ext_flash),
      .select_n_to_the_ext_flash_1             (select_n_to_the_ext_flash_1),
      .tb_fsm_address                          (tb_fsm_address),
      .tb_fsm_data                             (tb_fsm_data),
      .tb_fsm_readn                            (tb_fsm_readn),
      .tb_fsm_writen                           (tb_fsm_writen),
      .txd_from_the_uart                       (txd_from_the_uart),
      .txp_from_the_tse_mac                    (txp_from_the_tse_mac)
    );

  //default value specified in MODULE button_pio ptf port section
  assign in_port_to_the_button_pio = 7;

  //default value specified in MODULE dipsw_pio ptf port section
  assign in_port_to_the_dipsw_pio = 0;

  ext_flash the_ext_flash
    (
      .address  (tb_fsm_address[24 : 1]),
      .data     (tb_fsm_data),
      .read_n   (tb_fsm_readn),
      .select_n (select_n_to_the_ext_flash),
      .write_n  (tb_fsm_writen)
    );

  ext_flash_1 the_ext_flash_1
    (
      .address  (tb_fsm_address[24 : 1]),
      .data     (tb_fsm_data),
      .read_n   (tb_fsm_readn),
      .select_n (select_n_to_the_ext_flash_1),
      .write_n  (tb_fsm_writen)
    );

  tse_mac_loopback the_tse_mac_loopback
    (
      .ref_clk (ref_clk_to_the_tse_mac),
      .rxp     (rxp_to_the_tse_mac),
      .txp     (txp_from_the_tse_mac)
    );

  initial
    clkin_100 = 1'b0;
  always
    #5 clkin_100 <= ~clkin_100;
  
  initial 
    begin
      reset_n <= 0;
      #100 reset_n <= 1;
    end

endmodule


//synthesis translate_on